module edge_detection
(

);


endmodule