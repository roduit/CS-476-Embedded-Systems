module DMAController #(parameter [7:0] customId = 8'h00)
                    (input wire [31:0]  valueA,
                                        valueB,
                     output reg         status_register,
                     );



endmodule