--------------------------------------------------------------------------------
-- $RCSfile: $
--
-- DESC    : OpenRisk 1420 
--
-- AUTHOR  : Dr. Theo Kluter
--
-- CVS     : $Revision: $
--           $Date: $
--           $Author: $
--           $Source: $
--
--------------------------------------------------------------------------------
--
--  HISTORY :
--
--  $Log: 
--------------------------------------------------------------------------------

ARCHITECTURE platform_independent OF bios_rom IS

BEGIN

   TheRom : PROCESS( address )
   BEGIN
      CASE (address) IS
         WHEN "00000000000" => data <= X"EFBEADDE";
         WHEN "00000000001" => data <= X"00000015";
         WHEN "00000000010" => data <= X"21000000";
         WHEN "00000000011" => data <= X"00000015";
         WHEN "00000000100" => data <= X"1F000000";
         WHEN "00000000101" => data <= X"00000015";
         WHEN "00000000110" => data <= X"1D000000";
         WHEN "00000000111" => data <= X"00000015";
         WHEN "00000001000" => data <= X"1B000000";
         WHEN "00000001001" => data <= X"00000015";
         WHEN "00000001010" => data <= X"19000000";
         WHEN "00000001011" => data <= X"00000015";
         WHEN "00000001100" => data <= X"17000000";
         WHEN "00000001101" => data <= X"00000015";
         WHEN "00000001110" => data <= X"15000000";
         WHEN "00000001111" => data <= X"00000015";
         WHEN "00000010000" => data <= X"13000000";
         WHEN "00000010001" => data <= X"00000015";
         WHEN "00000010010" => data <= X"11000000";
         WHEN "00000010011" => data <= X"00000015";
         WHEN "00000010100" => data <= X"0F000000";
         WHEN "00000010101" => data <= X"00000015";
         WHEN "00000010110" => data <= X"0D000000";
         WHEN "00000010111" => data <= X"00000015";
         WHEN "00000011000" => data <= X"0B000000";
         WHEN "00000011001" => data <= X"00000015";
         WHEN "00000011010" => data <= X"09000000";
         WHEN "00000011011" => data <= X"00000015";
         WHEN "00000011100" => data <= X"00C02018";
         WHEN "00000011101" => data <= X"FC1F21A8";
         WHEN "00000011110" => data <= X"050060E0";
         WHEN "00000011111" => data <= X"FF020004";
         WHEN "00000100000" => data <= X"050080E0";
         WHEN "00000100010" => data <= X"00000015";
         WHEN "00000100011" => data <= X"84FF219C";
         WHEN "00000100100" => data <= X"001001D4";
         WHEN "00000100101" => data <= X"041801D4";
         WHEN "00000100110" => data <= X"082001D4";
         WHEN "00000100111" => data <= X"0C2801D4";
         WHEN "00000101000" => data <= X"103001D4";
         WHEN "00000101001" => data <= X"143801D4";
         WHEN "00000101010" => data <= X"184001D4";
         WHEN "00000101011" => data <= X"1C4801D4";
         WHEN "00000101100" => data <= X"205001D4";
         WHEN "00000101101" => data <= X"245801D4";
         WHEN "00000101110" => data <= X"286001D4";
         WHEN "00000101111" => data <= X"2C6801D4";
         WHEN "00000110000" => data <= X"307001D4";
         WHEN "00000110001" => data <= X"347801D4";
         WHEN "00000110010" => data <= X"388001D4";
         WHEN "00000110011" => data <= X"3C8801D4";
         WHEN "00000110100" => data <= X"409001D4";
         WHEN "00000110101" => data <= X"449801D4";
         WHEN "00000110110" => data <= X"48A001D4";
         WHEN "00000110111" => data <= X"4CA801D4";
         WHEN "00000111000" => data <= X"50B001D4";
         WHEN "00000111001" => data <= X"54B801D4";
         WHEN "00000111010" => data <= X"58C001D4";
         WHEN "00000111011" => data <= X"5CC801D4";
         WHEN "00000111100" => data <= X"60D001D4";
         WHEN "00000111101" => data <= X"64D801D4";
         WHEN "00000111110" => data <= X"68E001D4";
         WHEN "00000111111" => data <= X"6CE801D4";
         WHEN "00001000000" => data <= X"70F001D4";
         WHEN "00001000001" => data <= X"74F801D4";
         WHEN "00001000010" => data <= X"1200E0B7";
         WHEN "00001000011" => data <= X"0200FFBB";
         WHEN "00001000100" => data <= X"00F0C01B";
         WHEN "00001000101" => data <= X"AC01DEAB";
         WHEN "00001000110" => data <= X"00F8DEE3";
         WHEN "00001000111" => data <= X"0000FE87";
         WHEN "00001001000" => data <= X"00F80048";
         WHEN "00001001001" => data <= X"00000015";
         WHEN "00001001010" => data <= X"00004184";
         WHEN "00001001011" => data <= X"04006184";
         WHEN "00001001100" => data <= X"08008184";
         WHEN "00001001101" => data <= X"0C00A184";
         WHEN "00001001110" => data <= X"1000C184";
         WHEN "00001001111" => data <= X"1400E184";
         WHEN "00001010000" => data <= X"18000185";
         WHEN "00001010001" => data <= X"1C002185";
         WHEN "00001010010" => data <= X"20004185";
         WHEN "00001010011" => data <= X"24006185";
         WHEN "00001010100" => data <= X"28008185";
         WHEN "00001010101" => data <= X"2C00A185";
         WHEN "00001010110" => data <= X"3000C185";
         WHEN "00001010111" => data <= X"3400E185";
         WHEN "00001011000" => data <= X"38000186";
         WHEN "00001011001" => data <= X"3C002186";
         WHEN "00001011010" => data <= X"40004186";
         WHEN "00001011011" => data <= X"44006186";
         WHEN "00001011100" => data <= X"48008186";
         WHEN "00001011101" => data <= X"4C00A186";
         WHEN "00001011110" => data <= X"5000C186";
         WHEN "00001011111" => data <= X"5400E186";
         WHEN "00001100000" => data <= X"58000187";
         WHEN "00001100001" => data <= X"5C002187";
         WHEN "00001100010" => data <= X"60004187";
         WHEN "00001100011" => data <= X"64006187";
         WHEN "00001100100" => data <= X"68008187";
         WHEN "00001100101" => data <= X"6C00A187";
         WHEN "00001100110" => data <= X"7000C187";
         WHEN "00001100111" => data <= X"7400E187";
         WHEN "00001101000" => data <= X"7C00219C";
         WHEN "00001101001" => data <= X"00000024";
         WHEN "00001101010" => data <= X"00000015";
         WHEN "00001101011" => data <= X"700000F0";
         WHEN "00001101100" => data <= X"E40100F0";
         WHEN "00001101101" => data <= X"000200F0";
         WHEN "00001101110" => data <= X"1C0200F0";
         WHEN "00001101111" => data <= X"380200F0";
         WHEN "00001110000" => data <= X"540200F0";
         WHEN "00001110001" => data <= X"700200F0";
         WHEN "00001110010" => data <= X"8C0200F0";
         WHEN "00001110011" => data <= X"A80200F0";
         WHEN "00001110100" => data <= X"C40200F0";
         WHEN "00001110101" => data <= X"E00200F0";
         WHEN "00001110110" => data <= X"FC0200F0";
         WHEN "00001110111" => data <= X"340300F0";
         WHEN "00001111000" => data <= X"180300F0";
         WHEN "00001111001" => data <= X"00F0A018";
         WHEN "00001111010" => data <= X"00F08018";
         WHEN "00001111011" => data <= X"00F06018";
         WHEN "00001111100" => data <= X"E818A59C";
         WHEN "00001111101" => data <= X"B009849C";
         WHEN "00001111110" => data <= X"6A010000";
         WHEN "00001111111" => data <= X"180B639C";
         WHEN "00010000000" => data <= X"00F0A018";
         WHEN "00010000001" => data <= X"00F08018";
         WHEN "00010000010" => data <= X"00F06018";
         WHEN "00010000011" => data <= X"F418A59C";
         WHEN "00010000100" => data <= X"B009849C";
         WHEN "00010000101" => data <= X"63010000";
         WHEN "00010000110" => data <= X"180B639C";
         WHEN "00010000111" => data <= X"00F0A018";
         WHEN "00010001000" => data <= X"00F08018";
         WHEN "00010001001" => data <= X"00F06018";
         WHEN "00010001010" => data <= X"0519A59C";
         WHEN "00010001011" => data <= X"B009849C";
         WHEN "00010001100" => data <= X"5C010000";
         WHEN "00010001101" => data <= X"180B639C";
         WHEN "00010001110" => data <= X"00F0A018";
         WHEN "00010001111" => data <= X"00F08018";
         WHEN "00010010000" => data <= X"00F06018";
         WHEN "00010010001" => data <= X"1319A59C";
         WHEN "00010010010" => data <= X"B009849C";
         WHEN "00010010011" => data <= X"55010000";
         WHEN "00010010100" => data <= X"180B639C";
         WHEN "00010010101" => data <= X"00F0A018";
         WHEN "00010010110" => data <= X"00F08018";
         WHEN "00010010111" => data <= X"00F06018";
         WHEN "00010011000" => data <= X"1919A59C";
         WHEN "00010011001" => data <= X"B009849C";
         WHEN "00010011010" => data <= X"4E010000";
         WHEN "00010011011" => data <= X"180B639C";
         WHEN "00010011100" => data <= X"00F0A018";
         WHEN "00010011101" => data <= X"00F08018";
         WHEN "00010011110" => data <= X"00F06018";
         WHEN "00010011111" => data <= X"2219A59C";
         WHEN "00010100000" => data <= X"B009849C";
         WHEN "00010100001" => data <= X"47010000";
         WHEN "00010100010" => data <= X"180B639C";
         WHEN "00010100011" => data <= X"00F0A018";
         WHEN "00010100100" => data <= X"00F08018";
         WHEN "00010100101" => data <= X"00F06018";
         WHEN "00010100110" => data <= X"2819A59C";
         WHEN "00010100111" => data <= X"B009849C";
         WHEN "00010101000" => data <= X"40010000";
         WHEN "00010101001" => data <= X"180B639C";
         WHEN "00010101010" => data <= X"00F0A018";
         WHEN "00010101011" => data <= X"00F08018";
         WHEN "00010101100" => data <= X"00F06018";
         WHEN "00010101101" => data <= X"2E19A59C";
         WHEN "00010101110" => data <= X"B009849C";
         WHEN "00010101111" => data <= X"39010000";
         WHEN "00010110000" => data <= X"180B639C";
         WHEN "00010110001" => data <= X"00F0A018";
         WHEN "00010110010" => data <= X"00F08018";
         WHEN "00010110011" => data <= X"00F06018";
         WHEN "00010110100" => data <= X"3419A59C";
         WHEN "00010110101" => data <= X"B009849C";
         WHEN "00010110110" => data <= X"32010000";
         WHEN "00010110111" => data <= X"180B639C";
         WHEN "00010111000" => data <= X"00F0A018";
         WHEN "00010111001" => data <= X"00F08018";
         WHEN "00010111010" => data <= X"00F06018";
         WHEN "00010111011" => data <= X"3A19A59C";
         WHEN "00010111100" => data <= X"B009849C";
         WHEN "00010111101" => data <= X"2B010000";
         WHEN "00010111110" => data <= X"180B639C";
         WHEN "00010111111" => data <= X"00F0A018";
         WHEN "00011000000" => data <= X"00F08018";
         WHEN "00011000001" => data <= X"00F06018";
         WHEN "00011000010" => data <= X"4219A59C";
         WHEN "00011000011" => data <= X"B009849C";
         WHEN "00011000100" => data <= X"24010000";
         WHEN "00011000101" => data <= X"180B639C";
         WHEN "00011000110" => data <= X"00F0A018";
         WHEN "00011000111" => data <= X"00F08018";
         WHEN "00011001000" => data <= X"00F06018";
         WHEN "00011001001" => data <= X"4B19A59C";
         WHEN "00011001010" => data <= X"B009849C";
         WHEN "00011001011" => data <= X"1D010000";
         WHEN "00011001100" => data <= X"180B639C";
         WHEN "00011001101" => data <= X"00F0A018";
         WHEN "00011001110" => data <= X"00F08018";
         WHEN "00011001111" => data <= X"00F06018";
         WHEN "00011010000" => data <= X"5219A59C";
         WHEN "00011010001" => data <= X"B009849C";
         WHEN "00011010010" => data <= X"16010000";
         WHEN "00011010011" => data <= X"180B639C";
         WHEN "00011010100" => data <= X"0000601A";
         WHEN "00011010101" => data <= X"0700A0AA";
         WHEN "00011010110" => data <= X"02A83372";
         WHEN "00011010111" => data <= X"0000E01A";
         WHEN "00011011000" => data <= X"010031A6";
         WHEN "00011011001" => data <= X"00B831E4";
         WHEN "00011011010" => data <= X"FCFFFF13";
         WHEN "00011011011" => data <= X"00000015";
         WHEN "00011011100" => data <= X"00480044";
         WHEN "00011011101" => data <= X"00000015";
         WHEN "00011011110" => data <= X"00006019";
         WHEN "00011011111" => data <= X"02186B71";
         WHEN "00011100000" => data <= X"00480044";
         WHEN "00011100001" => data <= X"00000015";
         WHEN "00011100010" => data <= X"160020AA";
         WHEN "00011100011" => data <= X"02890370";
         WHEN "00011100100" => data <= X"020020AA";
         WHEN "00011100101" => data <= X"070060AA";
         WHEN "00011100110" => data <= X"02991170";
         WHEN "00011100111" => data <= X"EDFFFF03";
         WHEN "00011101000" => data <= X"00000015";
         WHEN "00011101001" => data <= X"DCFF219C";
         WHEN "00011101010" => data <= X"008001D4";
         WHEN "00011101011" => data <= X"049001D4";
         WHEN "00011101100" => data <= X"08A001D4";
         WHEN "00011101101" => data <= X"0CB001D4";
         WHEN "00011101110" => data <= X"10C001D4";
         WHEN "00011101111" => data <= X"14D001D4";
         WHEN "00011110000" => data <= X"18E001D4";
         WHEN "00011110001" => data <= X"1CF001D4";
         WHEN "00011110010" => data <= X"204801D4";
         WHEN "00011110011" => data <= X"0418C3E2";
         WHEN "00011110100" => data <= X"042044E2";
         WHEN "00011110101" => data <= X"0000001A";
         WHEN "00011110110" => data <= X"0000801A";
         WHEN "00011110111" => data <= X"160000AB";
         WHEN "00011111000" => data <= X"200040AB";
         WHEN "00011111001" => data <= X"010080AB";
         WHEN "00011111010" => data <= X"0700C0AB";
         WHEN "00011111011" => data <= X"009094E5";
         WHEN "00011111100" => data <= X"0C000010";
         WHEN "00011111101" => data <= X"20002185";
         WHEN "00011111110" => data <= X"00000186";
         WHEN "00011111111" => data <= X"04004186";
         WHEN "00100000000" => data <= X"08008186";
         WHEN "00100000001" => data <= X"0C00C186";
         WHEN "00100000010" => data <= X"10000187";
         WHEN "00100000011" => data <= X"14004187";
         WHEN "00100000100" => data <= X"18008187";
         WHEN "00100000101" => data <= X"1C00C187";
         WHEN "00100000110" => data <= X"00480044";
         WHEN "00100000111" => data <= X"2400219C";
         WHEN "00100001000" => data <= X"02C11070";
         WHEN "00100001001" => data <= X"180020AA";
         WHEN "00100001010" => data <= X"008076E2";
         WHEN "00100001011" => data <= X"0000B386";
         WHEN "00100001100" => data <= X"0102B572";
         WHEN "00100001101" => data <= X"02891570";
         WHEN "00100001110" => data <= X"0100319E";
         WHEN "00100001111" => data <= X"00D031E4";
         WHEN "00100010000" => data <= X"FBFFFF13";
         WHEN "00100010001" => data <= X"0400739E";
         WHEN "00100010010" => data <= X"02F11C70";
         WHEN "00100010011" => data <= X"C1FFFF07";
         WHEN "00100010100" => data <= X"0800949E";
         WHEN "00100010101" => data <= X"E6FFFF03";
         WHEN "00100010110" => data <= X"2000109E";
         WHEN "00100010111" => data <= X"B4FF219C";
         WHEN "00100011000" => data <= X"00F08018";
         WHEN "00100011001" => data <= X"2000A0A8";
         WHEN "00100011010" => data <= X"681E849C";
         WHEN "00100011011" => data <= X"0C00619C";
         WHEN "00100011100" => data <= X"2C8001D4";
         WHEN "00100011101" => data <= X"309001D4";
         WHEN "00100011110" => data <= X"38B001D4";
         WHEN "00100011111" => data <= X"3CC001D4";
         WHEN "00100100000" => data <= X"40D001D4";
         WHEN "00100100001" => data <= X"44E001D4";
         WHEN "00100100010" => data <= X"484801D4";
         WHEN "00100100011" => data <= X"34A001D4";
         WHEN "00100100100" => data <= X"A7010004";
         WHEN "00100100101" => data <= X"00F0401A";
         WHEN "00100100110" => data <= X"00F0001A";
         WHEN "00100100111" => data <= X"B009529E";
         WHEN "00100101000" => data <= X"180B109E";
         WHEN "00100101001" => data <= X"00F0A018";
         WHEN "00100101010" => data <= X"5919A59C";
         WHEN "00100101011" => data <= X"049092E0";
         WHEN "00100101100" => data <= X"BC000004";
         WHEN "00100101101" => data <= X"048070E0";
         WHEN "00100101110" => data <= X"1F00201A";
         WHEN "00100101111" => data <= X"00F0C01A";
         WHEN "00100110000" => data <= X"0000601A";
         WHEN "00100110001" => data <= X"00FC31AA";
         WHEN "00100110010" => data <= X"0004001B";
         WHEN "00100110011" => data <= X"FFFF40AF";
         WHEN "00100110100" => data <= X"8A19D69E";
         WHEN "00100110101" => data <= X"010080AB";
         WHEN "00100110110" => data <= X"0200A0AA";
         WHEN "00100110111" => data <= X"08A891E2";
         WHEN "00100111000" => data <= X"00C094E2";
         WHEN "00100111001" => data <= X"0000B486";
         WHEN "00100111010" => data <= X"00D015E4";
         WHEN "00100111011" => data <= X"1D000010";
         WHEN "00100111100" => data <= X"0100319E";
         WHEN "00100111101" => data <= X"0000201A";
         WHEN "00100111110" => data <= X"008813E4";
         WHEN "00100111111" => data <= X"10000010";
         WHEN "00101000000" => data <= X"04B0B6E0";
         WHEN "00101000001" => data <= X"00F0A018";
         WHEN "00101000010" => data <= X"7C19A59C";
         WHEN "00101000011" => data <= X"049092E0";
         WHEN "00101000100" => data <= X"048070E0";
         WHEN "00101000101" => data <= X"30004186";
         WHEN "00101000110" => data <= X"2C000186";
         WHEN "00101000111" => data <= X"34008186";
         WHEN "00101001000" => data <= X"3800C186";
         WHEN "00101001001" => data <= X"3C000187";
         WHEN "00101001010" => data <= X"40004187";
         WHEN "00101001011" => data <= X"44008187";
         WHEN "00101001100" => data <= X"48002185";
         WHEN "00101001101" => data <= X"9B000000";
         WHEN "00101001110" => data <= X"4C00219C";
         WHEN "00101001111" => data <= X"049092E0";
         WHEN "00101010000" => data <= X"98000004";
         WHEN "00101010001" => data <= X"048070E0";
         WHEN "00101010010" => data <= X"90FFFF07";
         WHEN "00101010011" => data <= X"04A074E0";
         WHEN "00101010100" => data <= X"1F00201A";
         WHEN "00101010101" => data <= X"04E07CE2";
         WHEN "00101010110" => data <= X"00FC31AA";
         WHEN "00101010111" => data <= X"0100319E";
         WHEN "00101011000" => data <= X"2000A01A";
         WHEN "00101011001" => data <= X"00A831E4";
         WHEN "00101011010" => data <= X"DDFFFF13";
         WHEN "00101011011" => data <= X"0200A0AA";
         WHEN "00101011100" => data <= X"00F0A018";
         WHEN "00101011101" => data <= X"A619A59C";
         WHEN "00101011110" => data <= X"049092E0";
         WHEN "00101011111" => data <= X"89000004";
         WHEN "00101100000" => data <= X"048070E0";
         WHEN "00101100001" => data <= X"0C00819E";
         WHEN "00101100010" => data <= X"04A074E2";
         WHEN "00101100011" => data <= X"180020AA";
         WHEN "00101100100" => data <= X"2000E0AA";
         WHEN "00101100101" => data <= X"0000B386";
         WHEN "00101100110" => data <= X"0102B572";
         WHEN "00101100111" => data <= X"02891570";
         WHEN "00101101000" => data <= X"0100319E";
         WHEN "00101101001" => data <= X"00B831E4";
         WHEN "00101101010" => data <= X"FBFFFF13";
         WHEN "00101101011" => data <= X"0400739E";
         WHEN "00101101100" => data <= X"7F00201A";
         WHEN "00101101101" => data <= X"00F031AA";
         WHEN "00101101110" => data <= X"160060AA";
         WHEN "00101101111" => data <= X"02991170";
         WHEN "00101110000" => data <= X"010020AA";
         WHEN "00101110001" => data <= X"070060AA";
         WHEN "00101110010" => data <= X"02991170";
         WHEN "00101110011" => data <= X"61FFFF07";
         WHEN "00101110100" => data <= X"00000015";
         WHEN "00101110101" => data <= X"00F0A018";
         WHEN "00101110110" => data <= X"C719A59C";
         WHEN "00101110111" => data <= X"049092E0";
         WHEN "00101111000" => data <= X"70000004";
         WHEN "00101111001" => data <= X"048070E0";
         WHEN "00101111010" => data <= X"7F04201A";
         WHEN "00101111011" => data <= X"00F031AA";
         WHEN "00101111100" => data <= X"0000601A";
         WHEN "00101111101" => data <= X"080020AB";
         WHEN "00101111110" => data <= X"0000B186";
         WHEN "00101111111" => data <= X"0000F486";
         WHEN "00110000000" => data <= X"00A817E4";
         WHEN "00110000001" => data <= X"14000010";
         WHEN "00110000010" => data <= X"0400319E";
         WHEN "00110000011" => data <= X"00F0A018";
         WHEN "00110000100" => data <= X"08B801D4";
         WHEN "00110000101" => data <= X"04A801D4";
         WHEN "00110000110" => data <= X"009801D4";
         WHEN "00110000111" => data <= X"049092E0";
         WHEN "00110001000" => data <= X"048070E0";
         WHEN "00110001001" => data <= X"5F000004";
         WHEN "00110001010" => data <= X"EC19A59C";
         WHEN "00110001011" => data <= X"48002185";
         WHEN "00110001100" => data <= X"2C000186";
         WHEN "00110001101" => data <= X"30004186";
         WHEN "00110001110" => data <= X"34008186";
         WHEN "00110001111" => data <= X"3800C186";
         WHEN "00110010000" => data <= X"3C000187";
         WHEN "00110010001" => data <= X"40004187";
         WHEN "00110010010" => data <= X"44008187";
         WHEN "00110010011" => data <= X"00480044";
         WHEN "00110010100" => data <= X"4C00219C";
         WHEN "00110010101" => data <= X"0100739E";
         WHEN "00110010110" => data <= X"00C833E4";
         WHEN "00110010111" => data <= X"E7FFFF13";
         WHEN "00110011000" => data <= X"0400949E";
         WHEN "00110011001" => data <= X"00F0A018";
         WHEN "00110011010" => data <= X"A9FFFF03";
         WHEN "00110011011" => data <= X"0C1AA59C";
         WHEN "00110011100" => data <= X"E8FF219C";
         WHEN "00110011101" => data <= X"008001D4";
         WHEN "00110011110" => data <= X"049001D4";
         WHEN "00110011111" => data <= X"08A001D4";
         WHEN "00110100000" => data <= X"0CB001D4";
         WHEN "00110100001" => data <= X"10C001D4";
         WHEN "00110100010" => data <= X"144801D4";
         WHEN "00110100011" => data <= X"041843E2";
         WHEN "00110100100" => data <= X"042084E2";
         WHEN "00110100101" => data <= X"1C0000AA";
         WHEN "00110100110" => data <= X"090000AB";
         WHEN "00110100111" => data <= X"FCFFC0AE";
         WHEN "00110101000" => data <= X"488074E0";
         WHEN "00110101001" => data <= X"0F0023A6";
         WHEN "00110101010" => data <= X"00C051E4";
         WHEN "00110101011" => data <= X"03000010";
         WHEN "00110101100" => data <= X"3700719C";
         WHEN "00110101101" => data <= X"3000719C";
         WHEN "00110101110" => data <= X"00900048";
         WHEN "00110101111" => data <= X"FCFF109E";
         WHEN "00110110000" => data <= X"00B030E4";
         WHEN "00110110001" => data <= X"F8FFFF13";
         WHEN "00110110010" => data <= X"488074E0";
         WHEN "00110110011" => data <= X"00000186";
         WHEN "00110110100" => data <= X"04004186";
         WHEN "00110110101" => data <= X"08008186";
         WHEN "00110110110" => data <= X"0C00C186";
         WHEN "00110110111" => data <= X"10000187";
         WHEN "00110111000" => data <= X"14002185";
         WHEN "00110111001" => data <= X"00480044";
         WHEN "00110111010" => data <= X"1800219C";
         WHEN "00110111011" => data <= X"E8FF219C";
         WHEN "00110111100" => data <= X"0C8001D4";
         WHEN "00110111101" => data <= X"109001D4";
         WHEN "00110111110" => data <= X"144801D4";
         WHEN "00110111111" => data <= X"041843E2";
         WHEN "00111000000" => data <= X"0000601A";
         WHEN "00111000001" => data <= X"0000001A";
         WHEN "00111000010" => data <= X"0A00A0AA";
         WHEN "00111000011" => data <= X"0AABE4E2";
         WHEN "00111000100" => data <= X"020020AA";
         WHEN "00111000101" => data <= X"088837E2";
         WHEN "00111000110" => data <= X"00B831E2";
         WHEN "00111000111" => data <= X"008831E2";
         WHEN "00111001000" => data <= X"028824E2";
         WHEN "00111001001" => data <= X"0200E19E";
         WHEN "00111001010" => data <= X"3000319E";
         WHEN "00111001011" => data <= X"0098F7E2";
         WHEN "00111001100" => data <= X"008817D8";
         WHEN "00111001101" => data <= X"0000201A";
         WHEN "00111001110" => data <= X"008813E4";
         WHEN "00111001111" => data <= X"04000010";
         WHEN "00111010000" => data <= X"008804E4";
         WHEN "00111010001" => data <= X"04000010";
         WHEN "00111010010" => data <= X"00000015";
         WHEN "00111010011" => data <= X"0100109E";
         WHEN "00111010100" => data <= X"FF0010A6";
         WHEN "00111010101" => data <= X"0100739E";
         WHEN "00111010110" => data <= X"00A833E4";
         WHEN "00111010111" => data <= X"ECFFFF13";
         WHEN "00111011000" => data <= X"0AAB84E0";
         WHEN "00111011001" => data <= X"0000201A";
         WHEN "00111011010" => data <= X"008830E4";
         WHEN "00111011011" => data <= X"07000010";
         WHEN "00111011100" => data <= X"FFFF109E";
         WHEN "00111011101" => data <= X"0C000186";
         WHEN "00111011110" => data <= X"10004186";
         WHEN "00111011111" => data <= X"14002185";
         WHEN "00111100000" => data <= X"00480044";
         WHEN "00111100001" => data <= X"1800219C";
         WHEN "00111100010" => data <= X"0200219E";
         WHEN "00111100011" => data <= X"008031E2";
         WHEN "00111100100" => data <= X"00900048";
         WHEN "00111100101" => data <= X"0000718C";
         WHEN "00111100110" => data <= X"F4FFFF03";
         WHEN "00111100111" => data <= X"0000201A";
         WHEN "00111101000" => data <= X"E0FF219C";
         WHEN "00111101001" => data <= X"008001D4";
         WHEN "00111101010" => data <= X"049001D4";
         WHEN "00111101011" => data <= X"08A001D4";
         WHEN "00111101100" => data <= X"0CB001D4";
         WHEN "00111101101" => data <= X"14D001D4";
         WHEN "00111101110" => data <= X"18E001D4";
         WHEN "00111101111" => data <= X"10C001D4";
         WHEN "00111110000" => data <= X"1C4801D4";
         WHEN "00111110001" => data <= X"041883E2";
         WHEN "00111110010" => data <= X"042004E2";
         WHEN "00111110011" => data <= X"042845E2";
         WHEN "00111110100" => data <= X"2000C19E";
         WHEN "00111110101" => data <= X"250040AB";
         WHEN "00111110110" => data <= X"630080AB";
         WHEN "00111110111" => data <= X"00007290";
         WHEN "00111111000" => data <= X"0000201A";
         WHEN "00111111001" => data <= X"008823E4";
         WHEN "00111111010" => data <= X"3B00000C";
         WHEN "00111111011" => data <= X"00D023E4";
         WHEN "00111111100" => data <= X"5A000010";
         WHEN "00111111101" => data <= X"FF0003A7";
         WHEN "00111111110" => data <= X"01003292";
         WHEN "00111111111" => data <= X"00E011E4";
         WHEN "01000000000" => data <= X"4D000010";
         WHEN "01000000001" => data <= X"00E051E5";
         WHEN "01000000010" => data <= X"1B000010";
         WHEN "01000000011" => data <= X"0000601A";
         WHEN "01000000100" => data <= X"009811E4";
         WHEN "01000000101" => data <= X"28000010";
         WHEN "01000000110" => data <= X"580060AA";
         WHEN "01000000111" => data <= X"009811E4";
         WHEN "01000001000" => data <= X"37000010";
         WHEN "01000001001" => data <= X"0400169F";
         WHEN "01000001010" => data <= X"00A00048";
         WHEN "01000001011" => data <= X"250060A8";
         WHEN "01000001100" => data <= X"0000201A";
         WHEN "01000001101" => data <= X"008810E4";
         WHEN "01000001110" => data <= X"04000010";
         WHEN "01000001111" => data <= X"00000015";
         WHEN "01000010000" => data <= X"00800048";
         WHEN "01000010001" => data <= X"250060A8";
         WHEN "01000010010" => data <= X"0100128F";
         WHEN "01000010011" => data <= X"00A00048";
         WHEN "01000010100" => data <= X"04C078E0";
         WHEN "01000010101" => data <= X"0000201A";
         WHEN "01000010110" => data <= X"008810E4";
         WHEN "01000010111" => data <= X"33000010";
         WHEN "01000011000" => data <= X"00000015";
         WHEN "01000011001" => data <= X"00800048";
         WHEN "01000011010" => data <= X"04C078E0";
         WHEN "01000011011" => data <= X"30000000";
         WHEN "01000011100" => data <= X"0100529E";
         WHEN "01000011101" => data <= X"640060AA";
         WHEN "01000011110" => data <= X"009811E4";
         WHEN "01000011111" => data <= X"EBFFFF0F";
         WHEN "01000100000" => data <= X"0400169F";
         WHEN "01000100001" => data <= X"04A074E0";
         WHEN "01000100010" => data <= X"0000D686";
         WHEN "01000100011" => data <= X"98FFFF07";
         WHEN "01000100100" => data <= X"04B096E0";
         WHEN "01000100101" => data <= X"0000201A";
         WHEN "01000100110" => data <= X"008810E4";
         WHEN "01000100111" => data <= X"22000010";
         WHEN "01000101000" => data <= X"04B096E0";
         WHEN "01000101001" => data <= X"92FFFF07";
         WHEN "01000101010" => data <= X"048070E0";
         WHEN "01000101011" => data <= X"1F000000";
         WHEN "01000101100" => data <= X"04C0D8E2";
         WHEN "01000101101" => data <= X"00A00048";
         WHEN "01000101110" => data <= X"04D07AE0";
         WHEN "01000101111" => data <= X"0000201A";
         WHEN "01000110000" => data <= X"008810E4";
         WHEN "01000110001" => data <= X"04000010";
         WHEN "01000110010" => data <= X"04D07AE0";
         WHEN "01000110011" => data <= X"00800048";
         WHEN "01000110100" => data <= X"00000015";
         WHEN "01000110101" => data <= X"00000186";
         WHEN "01000110110" => data <= X"04004186";
         WHEN "01000110111" => data <= X"08008186";
         WHEN "01000111000" => data <= X"0C00C186";
         WHEN "01000111001" => data <= X"10000187";
         WHEN "01000111010" => data <= X"14004187";
         WHEN "01000111011" => data <= X"18008187";
         WHEN "01000111100" => data <= X"1C002185";
         WHEN "01000111101" => data <= X"00480044";
         WHEN "01000111110" => data <= X"2000219C";
         WHEN "01000111111" => data <= X"04A074E0";
         WHEN "01001000000" => data <= X"0000D686";
         WHEN "01001000001" => data <= X"5BFFFF07";
         WHEN "01001000010" => data <= X"04B096E0";
         WHEN "01001000011" => data <= X"0000201A";
         WHEN "01001000100" => data <= X"008810E4";
         WHEN "01001000101" => data <= X"04000010";
         WHEN "01001000110" => data <= X"04B096E0";
         WHEN "01001000111" => data <= X"55FFFF07";
         WHEN "01001001000" => data <= X"048070E0";
         WHEN "01001001001" => data <= X"04C0D8E2";
         WHEN "01001001010" => data <= X"0100529E";
         WHEN "01001001011" => data <= X"ACFFFF03";
         WHEN "01001001100" => data <= X"0100529E";
         WHEN "01001001101" => data <= X"0300568E";
         WHEN "01001001110" => data <= X"00A00048";
         WHEN "01001001111" => data <= X"049072E0";
         WHEN "01001010000" => data <= X"0000201A";
         WHEN "01001010001" => data <= X"008810E4";
         WHEN "01001010010" => data <= X"E3FFFF13";
         WHEN "01001010011" => data <= X"049072E0";
         WHEN "01001010100" => data <= X"DFFFFF03";
         WHEN "01001010101" => data <= X"00000015";
         WHEN "01001010110" => data <= X"00A00048";
         WHEN "01001010111" => data <= X"04C078E0";
         WHEN "01001011000" => data <= X"0000201A";
         WHEN "01001011001" => data <= X"008810E4";
         WHEN "01001011010" => data <= X"F1FFFF13";
         WHEN "01001011011" => data <= X"00000015";
         WHEN "01001011100" => data <= X"00800048";
         WHEN "01001011101" => data <= X"04C078E0";
         WHEN "01001011110" => data <= X"99FFFF03";
         WHEN "01001011111" => data <= X"0100529E";
         WHEN "01001100000" => data <= X"0050201A";
         WHEN "01001100001" => data <= X"030071AA";
         WHEN "01001100010" => data <= X"83FFA0AE";
         WHEN "01001100011" => data <= X"00A813D8";
         WHEN "01001100100" => data <= X"1700A0AA";
         WHEN "01001100101" => data <= X"00A811D8";
         WHEN "01001100110" => data <= X"010031AA";
         WHEN "01001100111" => data <= X"000011D8";
         WHEN "01001101000" => data <= X"030020AA";
         WHEN "01001101001" => data <= X"008813D8";
         WHEN "01001101010" => data <= X"00480044";
         WHEN "01001101011" => data <= X"00000015";
         WHEN "01001101100" => data <= X"0050601A";
         WHEN "01001101101" => data <= X"FF0063A4";
         WHEN "01001101110" => data <= X"0500B3AA";
         WHEN "01001101111" => data <= X"0000358E";
         WHEN "01001110000" => data <= X"400031A6";
         WHEN "01001110001" => data <= X"0000E01A";
         WHEN "01001110010" => data <= X"00B811E4";
         WHEN "01001110011" => data <= X"05000010";
         WHEN "01001110100" => data <= X"00000015";
         WHEN "01001110101" => data <= X"001813D8";
         WHEN "01001110110" => data <= X"00480044";
         WHEN "01001110111" => data <= X"00000015";
         WHEN "01001111000" => data <= X"00000015";
         WHEN "01001111001" => data <= X"F6FFFF03";
         WHEN "01001111010" => data <= X"00000015";
         WHEN "01001111011" => data <= X"0050601A";
         WHEN "01001111100" => data <= X"0500B3AA";
         WHEN "01001111101" => data <= X"0000358E";
         WHEN "01001111110" => data <= X"010031A6";
         WHEN "01001111111" => data <= X"0000E01A";
         WHEN "01010000000" => data <= X"00B811E4";
         WHEN "01010000001" => data <= X"FCFFFF13";
         WHEN "01010000010" => data <= X"00000015";
         WHEN "01010000011" => data <= X"0000738D";
         WHEN "01010000100" => data <= X"00480044";
         WHEN "01010000101" => data <= X"00000015";
         WHEN "01010000110" => data <= X"F0FF219C";
         WHEN "01010000111" => data <= X"FF0063A4";
         WHEN "01010001000" => data <= X"008001D4";
         WHEN "01010001001" => data <= X"D0FF039E";
         WHEN "01010001010" => data <= X"FF0030A6";
         WHEN "01010001011" => data <= X"090060AA";
         WHEN "01010001100" => data <= X"049001D4";
         WHEN "01010001101" => data <= X"08A001D4";
         WHEN "01010001110" => data <= X"009851E4";
         WHEN "01010001111" => data <= X"0800000C";
         WHEN "01010010000" => data <= X"0C4801D4";
         WHEN "01010010001" => data <= X"BFFF239E";
         WHEN "01010010010" => data <= X"FF0031A6";
         WHEN "01010010011" => data <= X"050060AA";
         WHEN "01010010100" => data <= X"009851E4";
         WHEN "01010010101" => data <= X"18000010";
         WHEN "01010010110" => data <= X"C9FF039E";
         WHEN "01010010111" => data <= X"090040AA";
         WHEN "01010011000" => data <= X"050080AA";
         WHEN "01010011001" => data <= X"E2FFFF07";
         WHEN "01010011010" => data <= X"00000015";
         WHEN "01010011011" => data <= X"FF006BA5";
         WHEN "01010011100" => data <= X"D0FF2B9E";
         WHEN "01010011101" => data <= X"FF0071A6";
         WHEN "01010011110" => data <= X"009053E4";
         WHEN "01010011111" => data <= X"04000010";
         WHEN "01010100000" => data <= X"0400A0AA";
         WHEN "01010100001" => data <= X"08A810E2";
         WHEN "01010100010" => data <= X"008011E2";
         WHEN "01010100011" => data <= X"BFFF2B9E";
         WHEN "01010100100" => data <= X"FF0031A6";
         WHEN "01010100101" => data <= X"00A051E4";
         WHEN "01010100110" => data <= X"10000010";
         WHEN "01010100111" => data <= X"9FFF2B9E";
         WHEN "01010101000" => data <= X"040020AA";
         WHEN "01010101001" => data <= X"088810E2";
         WHEN "01010101010" => data <= X"C9FF6B9D";
         WHEN "01010101011" => data <= X"EEFFFF03";
         WHEN "01010101100" => data <= X"00800BE2";
         WHEN "01010101101" => data <= X"9FFF239E";
         WHEN "01010101110" => data <= X"FF0031A6";
         WHEN "01010101111" => data <= X"009851E4";
         WHEN "01010110000" => data <= X"04000010";
         WHEN "01010110001" => data <= X"00000015";
         WHEN "01010110010" => data <= X"E5FFFF03";
         WHEN "01010110011" => data <= X"A9FF039E";
         WHEN "01010110100" => data <= X"E3FFFF03";
         WHEN "01010110101" => data <= X"0000001A";
         WHEN "01010110110" => data <= X"FF0031A6";
         WHEN "01010110111" => data <= X"00A051E4";
         WHEN "01010111000" => data <= X"05000010";
         WHEN "01010111001" => data <= X"040020AA";
         WHEN "01010111010" => data <= X"088810E2";
         WHEN "01010111011" => data <= X"F0FFFF03";
         WHEN "01010111100" => data <= X"A9FF6B9D";
         WHEN "01010111101" => data <= X"0090B3E4";
         WHEN "01010111110" => data <= X"DBFFFF13";
         WHEN "01010111111" => data <= X"048070E1";
         WHEN "01011000000" => data <= X"04004186";
         WHEN "01011000001" => data <= X"00000186";
         WHEN "01011000010" => data <= X"08008186";
         WHEN "01011000011" => data <= X"0C002185";
         WHEN "01011000100" => data <= X"00480044";
         WHEN "01011000101" => data <= X"1000219C";
         WHEN "01011000110" => data <= X"FF0063A4";
         WHEN "01011000111" => data <= X"020020AA";
         WHEN "01011001000" => data <= X"00191170";
         WHEN "01011001001" => data <= X"00480044";
         WHEN "01011001010" => data <= X"00000015";
         WHEN "01011001011" => data <= X"041863E1";
         WHEN "01011001100" => data <= X"0000201A";
         WHEN "01011001101" => data <= X"002831E4";
         WHEN "01011001110" => data <= X"04000010";
         WHEN "01011001111" => data <= X"008864E2";
         WHEN "01011010000" => data <= X"00480044";
         WHEN "01011010001" => data <= X"00000015";
         WHEN "01011010010" => data <= X"0000B392";
         WHEN "01011010011" => data <= X"00886BE2";
         WHEN "01011010100" => data <= X"00A813D8";
         WHEN "01011010101" => data <= X"F8FFFF03";
         WHEN "01011010110" => data <= X"0100319E";
         WHEN "01011010111" => data <= X"E0FF219C";
         WHEN "01011011000" => data <= X"108001D4";
         WHEN "01011011001" => data <= X"149001D4";
         WHEN "01011011010" => data <= X"18A001D4";
         WHEN "01011011011" => data <= X"1C4801D4";
         WHEN "01011011100" => data <= X"030020AA";
         WHEN "01011011101" => data <= X"00011170";
         WHEN "01011011110" => data <= X"00F0801A";
         WHEN "01011011111" => data <= X"00F0401A";
         WHEN "01011100000" => data <= X"B009949E";
         WHEN "01011100001" => data <= X"180B529E";
         WHEN "01011100010" => data <= X"00F0A018";
         WHEN "01011100011" => data <= X"1F1AA59C";
         WHEN "01011100100" => data <= X"04A094E0";
         WHEN "01011100101" => data <= X"03FFFF07";
         WHEN "01011100110" => data <= X"049072E0";
         WHEN "01011100111" => data <= X"00F0A018";
         WHEN "01011101000" => data <= X"4E1AA59C";
         WHEN "01011101001" => data <= X"04A094E0";
         WHEN "01011101010" => data <= X"FEFEFF07";
         WHEN "01011101011" => data <= X"049072E0";
         WHEN "01011101100" => data <= X"00F0A018";
         WHEN "01011101101" => data <= X"711AA59C";
         WHEN "01011101110" => data <= X"04A094E0";
         WHEN "01011101111" => data <= X"F9FEFF07";
         WHEN "01011110000" => data <= X"049072E0";
         WHEN "01011110001" => data <= X"FF00201A";
         WHEN "01011110010" => data <= X"FFFF31AA";
         WHEN "01011110011" => data <= X"090000B6";
         WHEN "01011110100" => data <= X"0000A01A";
         WHEN "01011110101" => data <= X"038870E2";
         WHEN "01011110110" => data <= X"00A813E4";
         WHEN "01011110111" => data <= X"FCFFFF13";
         WHEN "01011111000" => data <= X"00F0A018";
         WHEN "01011111001" => data <= X"040020AA";
         WHEN "01011111010" => data <= X"488830E2";
         WHEN "01011111011" => data <= X"0F0031A6";
         WHEN "01011111100" => data <= X"048801D4";
         WHEN "01011111101" => data <= X"0F0030A6";
         WHEN "01011111110" => data <= X"008801D4";
         WHEN "01011111111" => data <= X"04A094E0";
         WHEN "01100000000" => data <= X"049072E0";
         WHEN "01100000001" => data <= X"E7FEFF07";
         WHEN "01100000010" => data <= X"9E1AA59C";
         WHEN "01100000011" => data <= X"0C0020AA";
         WHEN "01100000100" => data <= X"488830E2";
         WHEN "01100000101" => data <= X"0F0031A6";
         WHEN "01100000110" => data <= X"0C8801D4";
         WHEN "01100000111" => data <= X"100020AA";
         WHEN "01100001000" => data <= X"488830E2";
         WHEN "01100001001" => data <= X"0F0031A6";
         WHEN "01100001010" => data <= X"088801D4";
         WHEN "01100001011" => data <= X"140020AA";
         WHEN "01100001100" => data <= X"488830E2";
         WHEN "01100001101" => data <= X"0F0031A6";
         WHEN "01100001110" => data <= X"048801D4";
         WHEN "01100001111" => data <= X"180020AA";
         WHEN "01100010000" => data <= X"488810E2";
         WHEN "01100010001" => data <= X"0F0010A6";
         WHEN "01100010010" => data <= X"00F0A018";
         WHEN "01100010011" => data <= X"008001D4";
         WHEN "01100010100" => data <= X"04A094E0";
         WHEN "01100010101" => data <= X"049072E0";
         WHEN "01100010110" => data <= X"D2FEFF07";
         WHEN "01100010111" => data <= X"BC1AA59C";
         WHEN "01100011000" => data <= X"1C002185";
         WHEN "01100011001" => data <= X"10000186";
         WHEN "01100011010" => data <= X"14004186";
         WHEN "01100011011" => data <= X"18008186";
         WHEN "01100011100" => data <= X"00480044";
         WHEN "01100011101" => data <= X"2000219C";
         WHEN "01100011110" => data <= X"A4FC219C";
         WHEN "01100011111" => data <= X"307301D4";
         WHEN "01100100000" => data <= X"348301D4";
         WHEN "01100100001" => data <= X"389301D4";
         WHEN "01100100010" => data <= X"3CA301D4";
         WHEN "01100100011" => data <= X"40B301D4";
         WHEN "01100100100" => data <= X"44C301D4";
         WHEN "01100100101" => data <= X"48D301D4";
         WHEN "01100100110" => data <= X"4CE301D4";
         WHEN "01100100111" => data <= X"50F301D4";
         WHEN "01100101000" => data <= X"541301D4";
         WHEN "01100101001" => data <= X"584B01D4";
         WHEN "01100101010" => data <= X"00C0201A";
         WHEN "01100101011" => data <= X"068800C0";
         WHEN "01100101100" => data <= X"110020B6";
         WHEN "01100101101" => data <= X"2C8801D4";
         WHEN "01100101110" => data <= X"2C002186";
         WHEN "01100101111" => data <= X"100031AA";
         WHEN "01100110000" => data <= X"2C8801D4";
         WHEN "01100110001" => data <= X"2C002186";
         WHEN "01100110010" => data <= X"118800C0";
         WHEN "01100110011" => data <= X"2DFFFF07";
         WHEN "01100110100" => data <= X"010040AA";
         WHEN "01100110101" => data <= X"A2FFFF07";
         WHEN "01100110110" => data <= X"0000C01B";
         WHEN "01100110111" => data <= X"00F0201A";
         WHEN "01100111000" => data <= X"002031AA";
         WHEN "01100111001" => data <= X"0C8801D4";
         WHEN "01100111010" => data <= X"3F00201A";
         WHEN "01100111011" => data <= X"FFFF31AA";
         WHEN "01100111100" => data <= X"0000001B";
         WHEN "01100111101" => data <= X"0490D2E1";
         WHEN "01100111110" => data <= X"0000001A";
         WHEN "01100111111" => data <= X"188801D4";
         WHEN "01101000000" => data <= X"3BFFFF07";
         WHEN "01101000001" => data <= X"00000015";
         WHEN "01101000010" => data <= X"FF002BA6";
         WHEN "01101000011" => data <= X"270060AA";
         WHEN "01101000100" => data <= X"009811E4";
         WHEN "01101000101" => data <= X"87020010";
         WHEN "01101000110" => data <= X"04584BE3";
         WHEN "01101000111" => data <= X"009851E4";
         WHEN "01101001000" => data <= X"49000010";
         WHEN "01101001001" => data <= X"240060AA";
         WHEN "01101001010" => data <= X"009811E4";
         WHEN "01101001011" => data <= X"A1000010";
         WHEN "01101001100" => data <= X"009851E4";
         WHEN "01101001101" => data <= X"13000010";
         WHEN "01101001110" => data <= X"230060AA";
         WHEN "01101001111" => data <= X"009811E4";
         WHEN "01101010000" => data <= X"92000010";
         WHEN "01101010001" => data <= X"F6FF319E";
         WHEN "01101010010" => data <= X"FF0031A6";
         WHEN "01101010011" => data <= X"160060AA";
         WHEN "01101010100" => data <= X"009851E4";
         WHEN "01101010101" => data <= X"09000010";
         WHEN "01101010110" => data <= X"BFFF601A";
         WHEN "01101010111" => data <= X"F6FF73AA";
         WHEN "01101011000" => data <= X"888833E2";
         WHEN "01101011001" => data <= X"010031A6";
         WHEN "01101011010" => data <= X"0000601A";
         WHEN "01101011011" => data <= X"009831E4";
         WHEN "01101011100" => data <= X"E4FFFF0F";
         WHEN "01101011101" => data <= X"00000015";
         WHEN "01101011110" => data <= X"45000000";
         WHEN "01101011111" => data <= X"0000201A";
         WHEN "01101100000" => data <= X"260060AA";
         WHEN "01101100001" => data <= X"009811E4";
         WHEN "01101100010" => data <= X"4100000C";
         WHEN "01101100011" => data <= X"0000201A";
         WHEN "01101100100" => data <= X"17FFFF07";
         WHEN "01101100101" => data <= X"0000801B";
         WHEN "01101100110" => data <= X"00F0A018";
         WHEN "01101100111" => data <= X"00F08018";
         WHEN "01101101000" => data <= X"00F06018";
         WHEN "01101101001" => data <= X"DD1AA59C";
         WHEN "01101101010" => data <= X"B009849C";
         WHEN "01101101011" => data <= X"180B639C";
         WHEN "01101101100" => data <= X"7CFEFF07";
         WHEN "01101101101" => data <= X"FF004BA4";
         WHEN "01101101110" => data <= X"200040AB";
         WHEN "01101101111" => data <= X"00D002E4";
         WHEN "01101110000" => data <= X"1D000010";
         WHEN "01101110001" => data <= X"00E03CE2";
         WHEN "01101110010" => data <= X"00E031E2";
         WHEN "01101110011" => data <= X"3000619E";
         WHEN "01101110100" => data <= X"0088F3E2";
         WHEN "01101110101" => data <= X"0000A01A";
         WHEN "01101110110" => data <= X"0100B59E";
         WHEN "01101110111" => data <= X"001017D8";
         WHEN "01101111000" => data <= X"1C8801D4";
         WHEN "01101111001" => data <= X"14A801D4";
         WHEN "01101111010" => data <= X"01FFFF07";
         WHEN "01101111011" => data <= X"10B801D4";
         WHEN "01101111100" => data <= X"FF004BA4";
         WHEN "01101111101" => data <= X"00D022E4";
         WHEN "01101111110" => data <= X"1000E186";
         WHEN "01101111111" => data <= X"1400A186";
         WHEN "01110000000" => data <= X"0100F79E";
         WHEN "01110000001" => data <= X"F5FFFF13";
         WHEN "01110000010" => data <= X"1C002186";
         WHEN "01110000011" => data <= X"1003319E";
         WHEN "01110000100" => data <= X"2000619E";
         WHEN "01110000101" => data <= X"009831E2";
         WHEN "01110000110" => data <= X"00A831E2";
         WHEN "01110000111" => data <= X"0005F1DB";
         WHEN "01110001000" => data <= X"01009C9F";
         WHEN "01110001001" => data <= X"FF0020AA";
         WHEN "01110001010" => data <= X"0088BCE5";
         WHEN "01110001011" => data <= X"B5FFFF0F";
         WHEN "01110001100" => data <= X"00000015";
         WHEN "01110001101" => data <= X"EEFEFF07";
         WHEN "01110001110" => data <= X"00000015";
         WHEN "01110001111" => data <= X"E0FFFF03";
         WHEN "01110010000" => data <= X"FF004BA4";
         WHEN "01110010001" => data <= X"2D0060AA";
         WHEN "01110010010" => data <= X"009811E4";
         WHEN "01110010011" => data <= X"0B000010";
         WHEN "01110010100" => data <= X"009851E4";
         WHEN "01110010101" => data <= X"33000010";
         WHEN "01110010110" => data <= X"3D0060AA";
         WHEN "01110010111" => data <= X"2A0060AA";
         WHEN "01110011000" => data <= X"009811E4";
         WHEN "01110011001" => data <= X"62000010";
         WHEN "01110011010" => data <= X"2B0060AA";
         WHEN "01110011011" => data <= X"009811E4";
         WHEN "01110011100" => data <= X"0700000C";
         WHEN "01110011101" => data <= X"0000201A";
         WHEN "01110011110" => data <= X"DDFEFF07";
         WHEN "01110011111" => data <= X"00000015";
         WHEN "01110100000" => data <= X"180060AA";
         WHEN "01110100001" => data <= X"08982BE2";
         WHEN "01110100010" => data <= X"889831E2";
         WHEN "01110100011" => data <= X"180060AA";
         WHEN "01110100100" => data <= X"08987AE1";
         WHEN "01110100101" => data <= X"88986BE1";
         WHEN "01110100110" => data <= X"FFFF80AF";
         WHEN "01110100111" => data <= X"0000601A";
         WHEN "01110101000" => data <= X"FF00E0AA";
         WHEN "01110101001" => data <= X"0098B3E2";
         WHEN "01110101010" => data <= X"0098B5E2";
         WHEN "01110101011" => data <= X"2000219F";
         WHEN "01110101100" => data <= X"1003B59E";
         WHEN "01110101101" => data <= X"00C8B5E2";
         WHEN "01110101110" => data <= X"00FD3593";
         WHEN "01110101111" => data <= X"005839E4";
         WHEN "01110110000" => data <= X"08000010";
         WHEN "01110110001" => data <= X"00000015";
         WHEN "01110110010" => data <= X"01FDB592";
         WHEN "01110110011" => data <= X"008815E4";
         WHEN "01110110100" => data <= X"0400000C";
         WHEN "01110110101" => data <= X"00000015";
         WHEN "01110110110" => data <= X"049893E3";
         WHEN "01110110111" => data <= X"000160AA";
         WHEN "01110111000" => data <= X"0100739E";
         WHEN "01110111001" => data <= X"00B8B3E5";
         WHEN "01110111010" => data <= X"F0FFFF13";
         WHEN "01110111011" => data <= X"0098B3E2";
         WHEN "01110111100" => data <= X"0000201A";
         WHEN "01110111101" => data <= X"00887CE5";
         WHEN "01110111110" => data <= X"1B02000C";
         WHEN "01110111111" => data <= X"00F0A018";
         WHEN "01111000000" => data <= X"00F0401B";
         WHEN "01111000001" => data <= X"3A1E5A9F";
         WHEN "01111000010" => data <= X"0000201A";
         WHEN "01111000011" => data <= X"008832E4";
         WHEN "01111000100" => data <= X"18020010";
         WHEN "01111000101" => data <= X"00881EE4";
         WHEN "01111000110" => data <= X"7AFFFF03";
         WHEN "01111000111" => data <= X"010040AA";
         WHEN "01111001000" => data <= X"009811E4";
         WHEN "01111001001" => data <= X"D5FFFF13";
         WHEN "01111001010" => data <= X"400060AA";
         WHEN "01111001011" => data <= X"009811E4";
         WHEN "01111001100" => data <= X"D7FFFF0F";
         WHEN "01111001101" => data <= X"0000201A";
         WHEN "01111001110" => data <= X"B8FEFF07";
         WHEN "01111001111" => data <= X"200060A8";
         WHEN "01111010000" => data <= X"020020AA";
         WHEN "01111010001" => data <= X"00F0A018";
         WHEN "01111010010" => data <= X"00F06018";
         WHEN "01111010011" => data <= X"48888BE2";
         WHEN "01111010100" => data <= X"005801D4";
         WHEN "01111010101" => data <= X"18002186";
         WHEN "01111010110" => data <= X"F11AA59C";
         WHEN "01111010111" => data <= X"00008018";
         WHEN "01111011000" => data <= X"180B639C";
         WHEN "01111011001" => data <= X"038894E2";
         WHEN "01111011010" => data <= X"0EFEFF07";
         WHEN "01111011011" => data <= X"0458CBE2";
         WHEN "01111011100" => data <= X"0000201A";
         WHEN "01111011101" => data <= X"008814E4";
         WHEN "01111011110" => data <= X"62FFFF0F";
         WHEN "01111011111" => data <= X"0000C01B";
         WHEN "01111100000" => data <= X"60FFFF03";
         WHEN "01111100001" => data <= X"0000001B";
         WHEN "01111100010" => data <= X"00F0A018";
         WHEN "01111100011" => data <= X"CD1AA59C";
         WHEN "01111100100" => data <= X"00F08018";
         WHEN "01111100101" => data <= X"B009849C";
         WHEN "01111100110" => data <= X"00F06018";
         WHEN "01111100111" => data <= X"180B639C";
         WHEN "01111101000" => data <= X"00FEFF07";
         WHEN "01111101001" => data <= X"00000015";
         WHEN "01111101010" => data <= X"56FFFF03";
         WHEN "01111101011" => data <= X"00000015";
         WHEN "01111101100" => data <= X"ADDE201A";
         WHEN "01111101101" => data <= X"EFBE31AA";
         WHEN "01111101110" => data <= X"00007086";
         WHEN "01111101111" => data <= X"008813E4";
         WHEN "01111110000" => data <= X"05000010";
         WHEN "01111110001" => data <= X"0C002186";
         WHEN "01111110010" => data <= X"00F0A018";
         WHEN "01111110011" => data <= X"F1FFFF03";
         WHEN "01111110100" => data <= X"0F1BA59C";
         WHEN "01111110101" => data <= X"008830E4";
         WHEN "01111110110" => data <= X"93000010";
         WHEN "01111110111" => data <= X"010020AA";
         WHEN "01111111000" => data <= X"0F8880C3";
         WHEN "01111111001" => data <= X"47FFFF03";
         WHEN "01111111010" => data <= X"00000015";
         WHEN "01111111011" => data <= X"80FEFF07";
         WHEN "01111111100" => data <= X"00000015";
         WHEN "01111111101" => data <= X"FF006BA5";
         WHEN "01111111110" => data <= X"6D0020AA";
         WHEN "01111111111" => data <= X"00880BE4";
         WHEN "10000000000" => data <= X"6D010010";
         WHEN "10000000001" => data <= X"00884BE4";
         WHEN "10000000010" => data <= X"4F000010";
         WHEN "10000000011" => data <= X"730020AA";
         WHEN "10000000100" => data <= X"660020AA";
         WHEN "10000000101" => data <= X"00880BE4";
         WHEN "10000000110" => data <= X"13010010";
         WHEN "10000000111" => data <= X"00884BE4";
         WHEN "10000001000" => data <= X"32000010";
         WHEN "10000001001" => data <= X"680020AA";
         WHEN "10000001010" => data <= X"630020AA";
         WHEN "10000001011" => data <= X"00880BE4";
         WHEN "10000001100" => data <= X"CE000010";
         WHEN "10000001101" => data <= X"650020AA";
         WHEN "10000001110" => data <= X"00880BE4";
         WHEN "10000001111" => data <= X"31FFFF0F";
         WHEN "10000010000" => data <= X"00F0801B";
         WHEN "10000010001" => data <= X"00F0401B";
         WHEN "10000010010" => data <= X"B0099C9F";
         WHEN "10000010011" => data <= X"180B5A9F";
         WHEN "10000010100" => data <= X"00F0A018";
         WHEN "10000010101" => data <= X"041DA59C";
         WHEN "10000010110" => data <= X"04E09CE0";
         WHEN "10000010111" => data <= X"D1FDFF07";
         WHEN "10000011000" => data <= X"04D07AE0";
         WHEN "10000011001" => data <= X"00F0A018";
         WHEN "10000011010" => data <= X"00044018";
         WHEN "10000011011" => data <= X"FFFFA0AE";
         WHEN "10000011100" => data <= X"00FCE01A";
         WHEN "10000011101" => data <= X"AE1CA59C";
         WHEN "10000011110" => data <= X"0005601A";
         WHEN "10000011111" => data <= X"00002286";
         WHEN "10000100000" => data <= X"00A811E4";
         WHEN "10000100001" => data <= X"12000010";
         WHEN "10000100010" => data <= X"00B822E2";
         WHEN "10000100011" => data <= X"008801D4";
         WHEN "10000100100" => data <= X"04E09CE0";
         WHEN "10000100101" => data <= X"04D07AE0";
         WHEN "10000100110" => data <= X"249801D4";
         WHEN "10000100111" => data <= X"20A801D4";
         WHEN "10000101000" => data <= X"1CB801D4";
         WHEN "10000101001" => data <= X"102801D4";
         WHEN "10000101010" => data <= X"BEFDFF07";
         WHEN "10000101011" => data <= X"148801D4";
         WHEN "10000101100" => data <= X"14002186";
         WHEN "10000101101" => data <= X"B5FCFF07";
         WHEN "10000101110" => data <= X"048871E0";
         WHEN "10000101111" => data <= X"24006186";
         WHEN "10000110000" => data <= X"2000A186";
         WHEN "10000110001" => data <= X"1C00E186";
         WHEN "10000110010" => data <= X"1000A184";
         WHEN "10000110011" => data <= X"0400429C";
         WHEN "10000110100" => data <= X"009822E4";
         WHEN "10000110101" => data <= X"EAFFFF13";
         WHEN "10000110110" => data <= X"00000015";
         WHEN "10000110111" => data <= X"00F0A018";
         WHEN "10000111000" => data <= X"EF000000";
         WHEN "10000111001" => data <= X"221DA59C";
         WHEN "10000111010" => data <= X"00880BE4";
         WHEN "10000111011" => data <= X"38000010";
         WHEN "10000111100" => data <= X"690020AA";
         WHEN "10000111101" => data <= X"00880BE4";
         WHEN "10000111110" => data <= X"02FFFF0F";
         WHEN "10000111111" => data <= X"ADDE201A";
         WHEN "10001000000" => data <= X"EFBE31AA";
         WHEN "10001000001" => data <= X"00007086";
         WHEN "10001000010" => data <= X"00F08018";
         WHEN "10001000011" => data <= X"008813E4";
         WHEN "10001000100" => data <= X"00F06018";
         WHEN "10001000101" => data <= X"04003086";
         WHEN "10001000110" => data <= X"B009849C";
         WHEN "10001000111" => data <= X"6B000010";
         WHEN "10001001000" => data <= X"180B639C";
         WHEN "10001001001" => data <= X"00F0A018";
         WHEN "10001001010" => data <= X"048801D4";
         WHEN "10001001011" => data <= X"000001D4";
         WHEN "10001001100" => data <= X"851BA59C";
         WHEN "10001001101" => data <= X"9BFDFF07";
         WHEN "10001001110" => data <= X"00000015";
         WHEN "10001001111" => data <= X"F1FEFF03";
         WHEN "10001010000" => data <= X"00000015";
         WHEN "10001010001" => data <= X"00880BE4";
         WHEN "10001010010" => data <= X"2B000010";
         WHEN "10001010011" => data <= X"00884BE4";
         WHEN "10001010100" => data <= X"11000010";
         WHEN "10001010101" => data <= X"740020AA";
         WHEN "10001010110" => data <= X"700020AA";
         WHEN "10001010111" => data <= X"00880BE4";
         WHEN "10001011000" => data <= X"51000010";
         WHEN "10001011001" => data <= X"720020AA";
         WHEN "10001011010" => data <= X"00880BE4";
         WHEN "10001011011" => data <= X"E5FEFF0F";
         WHEN "10001011100" => data <= X"ADDE201A";
         WHEN "10001011101" => data <= X"0004A01A";
         WHEN "10001011110" => data <= X"EFBE31AA";
         WHEN "10001011111" => data <= X"00007586";
         WHEN "10001100000" => data <= X"008813E4";
         WHEN "10001100001" => data <= X"20000010";
         WHEN "10001100010" => data <= X"00F0A018";
         WHEN "10001100011" => data <= X"81FFFF03";
         WHEN "10001100100" => data <= X"3F1BA59C";
         WHEN "10001100101" => data <= X"00880BE4";
         WHEN "10001100110" => data <= X"55000010";
         WHEN "10001100111" => data <= X"760020AA";
         WHEN "10001101000" => data <= X"00880BE4";
         WHEN "10001101001" => data <= X"D7FEFF0F";
         WHEN "10001101010" => data <= X"00F0A018";
         WHEN "10001101011" => data <= X"00F08018";
         WHEN "10001101100" => data <= X"00F06018";
         WHEN "10001101101" => data <= X"701BA59C";
         WHEN "10001101110" => data <= X"B009849C";
         WHEN "10001101111" => data <= X"79FDFF07";
         WHEN "10001110000" => data <= X"180B639C";
         WHEN "10001110001" => data <= X"CFFEFF03";
         WHEN "10001110010" => data <= X"0000C019";
         WHEN "10001110011" => data <= X"00F0A018";
         WHEN "10001110100" => data <= X"00F06018";
         WHEN "10001110101" => data <= X"3A1DA59C";
         WHEN "10001110110" => data <= X"00008018";
         WHEN "10001110111" => data <= X"71FDFF07";
         WHEN "10001111000" => data <= X"B009639C";
         WHEN "10001111001" => data <= X"5EFEFF07";
         WHEN "10001111010" => data <= X"00000015";
         WHEN "10001111011" => data <= X"C5FEFF03";
         WHEN "10001111100" => data <= X"00000015";
         WHEN "10001111101" => data <= X"9AFCFF07";
         WHEN "10001111110" => data <= X"00000015";
         WHEN "10001111111" => data <= X"C1FEFF03";
         WHEN "10010000000" => data <= X"00000015";
         WHEN "10010000001" => data <= X"040035AA";
         WHEN "10010000010" => data <= X"00007186";
         WHEN "10010000011" => data <= X"020020AA";
         WHEN "10010000100" => data <= X"088873E2";
         WHEN "10010000101" => data <= X"0000201A";
         WHEN "10010000110" => data <= X"009831E4";
         WHEN "10010000111" => data <= X"1D000010";
         WHEN "10010001000" => data <= X"0088F5E2";
         WHEN "10010001001" => data <= X"110020B6";
         WHEN "10010001010" => data <= X"FFBF60AE";
         WHEN "10010001011" => data <= X"2C8801D4";
         WHEN "10010001100" => data <= X"2C002186";
         WHEN "10010001101" => data <= X"039831E2";
         WHEN "10010001110" => data <= X"2C8801D4";
         WHEN "10010001111" => data <= X"2C002186";
         WHEN "10010010000" => data <= X"118800C0";
         WHEN "10010010001" => data <= X"E7BF60AE";
         WHEN "10010010010" => data <= X"2C002186";
         WHEN "10010010011" => data <= X"039831E2";
         WHEN "10010010100" => data <= X"2C8801D4";
         WHEN "10010010101" => data <= X"0D0040AB";
         WHEN "10010010110" => data <= X"00E05AB7";
         WHEN "10010010111" => data <= X"00F0A018";
         WHEN "10010011000" => data <= X"00F08018";
         WHEN "10010011001" => data <= X"00F06018";
         WHEN "10010011010" => data <= X"2A1BA59C";
         WHEN "10010011011" => data <= X"B009849C";
         WHEN "10010011100" => data <= X"4CFDFF07";
         WHEN "10010011101" => data <= X"180B639C";
         WHEN "10010011110" => data <= X"04D050E3";
         WHEN "10010011111" => data <= X"2C002186";
         WHEN "10010100000" => data <= X"00D00044";
         WHEN "10010100001" => data <= X"118800C0";
         WHEN "10010100010" => data <= X"9EFEFF03";
         WHEN "10010100011" => data <= X"00000015";
         WHEN "10010100100" => data <= X"0000F786";
         WHEN "10010100101" => data <= X"0400319E";
         WHEN "10010100110" => data <= X"FCBFF1D7";
         WHEN "10010100111" => data <= X"E0FFFF03";
         WHEN "10010101000" => data <= X"009831E4";
         WHEN "10010101001" => data <= X"00F0A018";
         WHEN "10010101010" => data <= X"00F08018";
         WHEN "10010101011" => data <= X"00F06018";
         WHEN "10010101100" => data <= X"5C1BA59C";
         WHEN "10010101101" => data <= X"B009849C";
         WHEN "10010101110" => data <= X"3AFDFF07";
         WHEN "10010101111" => data <= X"180B639C";
         WHEN "10010110000" => data <= X"90FEFF03";
         WHEN "10010110001" => data <= X"0100C0A9";
         WHEN "10010110010" => data <= X"020060AA";
         WHEN "10010110011" => data <= X"089831E2";
         WHEN "10010110100" => data <= X"048031E2";
         WHEN "10010110101" => data <= X"FFFF319E";
         WHEN "10010110110" => data <= X"00F0A018";
         WHEN "10010110111" => data <= X"048801D4";
         WHEN "10010111000" => data <= X"008001D4";
         WHEN "10010111001" => data <= X"94FFFF03";
         WHEN "10010111010" => data <= X"991BA59C";
         WHEN "10010111011" => data <= X"0000201A";
         WHEN "10010111100" => data <= X"00F08018";
         WHEN "10010111101" => data <= X"00F06018";
         WHEN "10010111110" => data <= X"008830E4";
         WHEN "10010111111" => data <= X"B009849C";
         WHEN "10011000000" => data <= X"09000010";
         WHEN "10011000001" => data <= X"180B639C";
         WHEN "10011000010" => data <= X"00F0A018";
         WHEN "10011000011" => data <= X"BB1BA59C";
         WHEN "10011000100" => data <= X"24FDFF07";
         WHEN "10011000101" => data <= X"00F0001A";
         WHEN "10011000110" => data <= X"0000001B";
         WHEN "10011000111" => data <= X"79FEFF03";
         WHEN "10011001000" => data <= X"002010AA";
         WHEN "10011001001" => data <= X"00F0201A";
         WHEN "10011001010" => data <= X"002031AA";
         WHEN "10011001011" => data <= X"008830E4";
         WHEN "10011001100" => data <= X"08000010";
         WHEN "10011001101" => data <= X"00000015";
         WHEN "10011001110" => data <= X"00F0A018";
         WHEN "10011001111" => data <= X"19FDFF07";
         WHEN "10011010000" => data <= X"D21BA59C";
         WHEN "10011010001" => data <= X"0000001B";
         WHEN "10011010010" => data <= X"6EFEFF03";
         WHEN "10011010011" => data <= X"0004001A";
         WHEN "10011010100" => data <= X"00F0A018";
         WHEN "10011010101" => data <= X"13FDFF07";
         WHEN "10011010110" => data <= X"E51BA59C";
         WHEN "10011010111" => data <= X"0000001B";
         WHEN "10011011000" => data <= X"68FEFF03";
         WHEN "10011011001" => data <= X"0000001A";
         WHEN "10011011010" => data <= X"00F0201A";
         WHEN "10011011011" => data <= X"002031AA";
         WHEN "10011011100" => data <= X"008810E4";
         WHEN "10011011101" => data <= X"05000010";
         WHEN "10011011110" => data <= X"0004201A";
         WHEN "10011011111" => data <= X"008830E4";
         WHEN "10011100000" => data <= X"05000010";
         WHEN "10011100001" => data <= X"ADDE201A";
         WHEN "10011100010" => data <= X"00F0A018";
         WHEN "10011100011" => data <= X"01FFFF03";
         WHEN "10011100100" => data <= X"F81BA59C";
         WHEN "10011100101" => data <= X"EFBE31AA";
         WHEN "10011100110" => data <= X"00007086";
         WHEN "10011100111" => data <= X"008813E4";
         WHEN "10011101000" => data <= X"05000010";
         WHEN "10011101001" => data <= X"3F00201A";
         WHEN "10011101010" => data <= X"00F0A018";
         WHEN "10011101011" => data <= X"F9FEFF03";
         WHEN "10011101100" => data <= X"1A1CA59C";
         WHEN "10011101101" => data <= X"FFFF31AA";
         WHEN "10011101110" => data <= X"04007086";
         WHEN "10011101111" => data <= X"0088B3E4";
         WHEN "10011110000" => data <= X"21000010";
         WHEN "10011110001" => data <= X"00F0A018";
         WHEN "10011110010" => data <= X"F2FEFF03";
         WHEN "10011110011" => data <= X"371CA59C";
         WHEN "10011110100" => data <= X"0088BAE2";
         WHEN "10011110101" => data <= X"00007587";
         WHEN "10011110110" => data <= X"00003A87";
         WHEN "10011110111" => data <= X"00C81BE4";
         WHEN "10011111000" => data <= X"10000010";
         WHEN "10011111001" => data <= X"04883AE2";
         WHEN "10011111010" => data <= X"00F06018";
         WHEN "10011111011" => data <= X"0000B586";
         WHEN "10011111100" => data <= X"0410A2E0";
         WHEN "10011111101" => data <= X"00003A87";
         WHEN "10011111110" => data <= X"04E09CE0";
         WHEN "10011111111" => data <= X"08C801D4";
         WHEN "10100000000" => data <= X"04A801D4";
         WHEN "10100000001" => data <= X"008801D4";
         WHEN "10100000010" => data <= X"180B639C";
         WHEN "10100000011" => data <= X"14B801D4";
         WHEN "10100000100" => data <= X"E4FCFF07";
         WHEN "10100000101" => data <= X"109801D4";
         WHEN "10100000110" => data <= X"1400E186";
         WHEN "10100000111" => data <= X"10006186";
         WHEN "10100001000" => data <= X"0100739E";
         WHEN "10100001001" => data <= X"04005A9F";
         WHEN "10100001010" => data <= X"00003786";
         WHEN "10100001011" => data <= X"009851E4";
         WHEN "10100001100" => data <= X"E8FFFF13";
         WHEN "10100001101" => data <= X"0004201A";
         WHEN "10100001110" => data <= X"00F0A018";
         WHEN "10100001111" => data <= X"D5FEFF03";
         WHEN "10100010000" => data <= X"7D1CA59C";
         WHEN "10100010001" => data <= X"00F04018";
         WHEN "10100010010" => data <= X"00F0801B";
         WHEN "10100010011" => data <= X"0000401B";
         WHEN "10100010100" => data <= X"0000601A";
         WHEN "10100010101" => data <= X"0400E0AA";
         WHEN "10100010110" => data <= X"571C429C";
         WHEN "10100010111" => data <= X"F3FFFF03";
         WHEN "10100011000" => data <= X"B0099C9F";
         WHEN "10100011001" => data <= X"00F0201A";
         WHEN "10100011010" => data <= X"002031AA";
         WHEN "10100011011" => data <= X"00F0801B";
         WHEN "10100011100" => data <= X"00F0401B";
         WHEN "10100011101" => data <= X"008810E4";
         WHEN "10100011110" => data <= X"B0099C9F";
         WHEN "10100011111" => data <= X"06000010";
         WHEN "10100100000" => data <= X"180B5A9F";
         WHEN "10100100001" => data <= X"0004201A";
         WHEN "10100100010" => data <= X"008830E4";
         WHEN "10100100011" => data <= X"07000010";
         WHEN "10100100100" => data <= X"ADDE201A";
         WHEN "10100100101" => data <= X"00F0A018";
         WHEN "10100100110" => data <= X"F81BA59C";
         WHEN "10100100111" => data <= X"04E09CE0";
         WHEN "10100101000" => data <= X"C0FEFF03";
         WHEN "10100101001" => data <= X"04D07AE0";
         WHEN "10100101010" => data <= X"EFBE31AA";
         WHEN "10100101011" => data <= X"00007086";
         WHEN "10100101100" => data <= X"008813E4";
         WHEN "10100101101" => data <= X"05000010";
         WHEN "10100101110" => data <= X"3F00201A";
         WHEN "10100101111" => data <= X"00F0A018";
         WHEN "10100110000" => data <= X"F7FFFF03";
         WHEN "10100110001" => data <= X"1A1CA59C";
         WHEN "10100110010" => data <= X"FFFF31AA";
         WHEN "10100110011" => data <= X"04007086";
         WHEN "10100110100" => data <= X"0088B3E4";
         WHEN "10100110101" => data <= X"04000010";
         WHEN "10100110110" => data <= X"00F0A018";
         WHEN "10100110111" => data <= X"F0FFFF03";
         WHEN "10100111000" => data <= X"371CA59C";
         WHEN "10100111001" => data <= X"00F0A018";
         WHEN "10100111010" => data <= X"8B1CA59C";
         WHEN "10100111011" => data <= X"04E09CE0";
         WHEN "10100111100" => data <= X"ACFCFF07";
         WHEN "10100111101" => data <= X"04D07AE0";
         WHEN "10100111110" => data <= X"00F0A018";
         WHEN "10100111111" => data <= X"0004201A";
         WHEN "10101000000" => data <= X"0000601A";
         WHEN "10101000001" => data <= X"040040A8";
         WHEN "10101000010" => data <= X"FFFFE0AE";
         WHEN "10101000011" => data <= X"00FC201B";
         WHEN "10101000100" => data <= X"AE1CA59C";
         WHEN "10101000101" => data <= X"0000A286";
         WHEN "10101000110" => data <= X"009855E4";
         WHEN "10101000111" => data <= X"0D000010";
         WHEN "10101001000" => data <= X"04E09CE0";
         WHEN "10101001001" => data <= X"00F0A018";
         WHEN "10101001010" => data <= X"D51CA59C";
         WHEN "10101001011" => data <= X"9DFCFF07";
         WHEN "10101001100" => data <= X"04D07AE0";
         WHEN "10101001101" => data <= X"00006018";
         WHEN "10101001110" => data <= X"00008284";
         WHEN "10101001111" => data <= X"9AFBFF07";
         WHEN "10101010000" => data <= X"00000015";
         WHEN "10101010001" => data <= X"00F0A018";
         WHEN "10101010010" => data <= X"D5FFFF03";
         WHEN "10101010011" => data <= X"EE1CA59C";
         WHEN "10101010100" => data <= X"0000B186";
         WHEN "10101010101" => data <= X"00B815E4";
         WHEN "10101010110" => data <= X"14000010";
         WHEN "10101010111" => data <= X"00C8B1E2";
         WHEN "10101011000" => data <= X"00A801D4";
         WHEN "10101011001" => data <= X"04E09CE0";
         WHEN "10101011010" => data <= X"04D07AE0";
         WHEN "10101011011" => data <= X"28B801D4";
         WHEN "10101011100" => data <= X"249801D4";
         WHEN "10101011101" => data <= X"20C801D4";
         WHEN "10101011110" => data <= X"1C8801D4";
         WHEN "10101011111" => data <= X"102801D4";
         WHEN "10101100000" => data <= X"88FCFF07";
         WHEN "10101100001" => data <= X"14A801D4";
         WHEN "10101100010" => data <= X"1400A186";
         WHEN "10101100011" => data <= X"7FFBFF07";
         WHEN "10101100100" => data <= X"04A875E0";
         WHEN "10101100101" => data <= X"2800E186";
         WHEN "10101100110" => data <= X"24006186";
         WHEN "10101100111" => data <= X"20002187";
         WHEN "10101101000" => data <= X"1C002186";
         WHEN "10101101001" => data <= X"1000A184";
         WHEN "10101101010" => data <= X"0100739E";
         WHEN "10101101011" => data <= X"DAFFFF03";
         WHEN "10101101100" => data <= X"0400319E";
         WHEN "10101101101" => data <= X"00F0401B";
         WHEN "10101101110" => data <= X"00F0001B";
         WHEN "10101101111" => data <= X"B0095A9F";
         WHEN "10101110000" => data <= X"180B189F";
         WHEN "10101110001" => data <= X"00F0A018";
         WHEN "10101110010" => data <= X"3D1DA59C";
         WHEN "10101110011" => data <= X"04D09AE0";
         WHEN "10101110100" => data <= X"74FCFF07";
         WHEN "10101110101" => data <= X"04C078E0";
         WHEN "10101110110" => data <= X"00F0201A";
         WHEN "10101110111" => data <= X"5F1D319E";
         WHEN "10101111000" => data <= X"108801D4";
         WHEN "10101111001" => data <= X"00F0201A";
         WHEN "10101111010" => data <= X"791D319E";
         WHEN "10101111011" => data <= X"0000801B";
         WHEN "10101111100" => data <= X"148801D4";
         WHEN "10101111101" => data <= X"04D09AE0";
         WHEN "10101111110" => data <= X"04C078E0";
         WHEN "10101111111" => data <= X"69FCFF07";
         WHEN "10110000000" => data <= X"1000A184";
         WHEN "10110000001" => data <= X"0000201A";
         WHEN "10110000010" => data <= X"0002601A";
         WHEN "10110000011" => data <= X"0200A0AA";
         WHEN "10110000100" => data <= X"00A81CE4";
         WHEN "10110000101" => data <= X"03000010";
         WHEN "10110000110" => data <= X"00000015";
         WHEN "10110000111" => data <= X"0100F172";
         WHEN "10110001000" => data <= X"008811D4";
         WHEN "10110001001" => data <= X"0400319E";
         WHEN "10110001010" => data <= X"009831E4";
         WHEN "10110001011" => data <= X"F9FFFF13";
         WHEN "10110001100" => data <= X"0200A0AA";
         WHEN "10110001101" => data <= X"00F0A018";
         WHEN "10110001110" => data <= X"6B1DA59C";
         WHEN "10110001111" => data <= X"04D09AE0";
         WHEN "10110010000" => data <= X"58FCFF07";
         WHEN "10110010001" => data <= X"04C078E0";
         WHEN "10110010010" => data <= X"0000201A";
         WHEN "10110010011" => data <= X"00004018";
         WHEN "10110010100" => data <= X"1D0020AB";
         WHEN "10110010101" => data <= X"0002E01A";
         WHEN "10110010110" => data <= X"020060AA";
         WHEN "10110010111" => data <= X"00981CE4";
         WHEN "10110011000" => data <= X"03000010";
         WHEN "10110011001" => data <= X"00000015";
         WHEN "10110011010" => data <= X"01007173";
         WHEN "10110011011" => data <= X"00007187";
         WHEN "10110011100" => data <= X"00881BE4";
         WHEN "10110011101" => data <= X"13000010";
         WHEN "10110011110" => data <= X"00C842E4";
         WHEN "10110011111" => data <= X"10000010";
         WHEN "10110100000" => data <= X"00000015";
         WHEN "10110100001" => data <= X"00007187";
         WHEN "10110100010" => data <= X"04D09AE0";
         WHEN "10110100011" => data <= X"088801D4";
         WHEN "10110100100" => data <= X"008801D4";
         WHEN "10110100101" => data <= X"04D801D4";
         WHEN "10110100110" => data <= X"04C078E0";
         WHEN "10110100111" => data <= X"24C801D4";
         WHEN "10110101000" => data <= X"20B801D4";
         WHEN "10110101001" => data <= X"1C8801D4";
         WHEN "10110101010" => data <= X"3EFCFF07";
         WHEN "10110101011" => data <= X"1400A184";
         WHEN "10110101100" => data <= X"24002187";
         WHEN "10110101101" => data <= X"2000E186";
         WHEN "10110101110" => data <= X"1C002186";
         WHEN "10110101111" => data <= X"0100429C";
         WHEN "10110110000" => data <= X"0400319E";
         WHEN "10110110001" => data <= X"00B831E4";
         WHEN "10110110010" => data <= X"E5FFFF13";
         WHEN "10110110011" => data <= X"020060AA";
         WHEN "10110110100" => data <= X"0000201A";
         WHEN "10110110101" => data <= X"008802E4";
         WHEN "10110110110" => data <= X"10000010";
         WHEN "10110110111" => data <= X"030020AA";
         WHEN "10110111000" => data <= X"00F0A018";
         WHEN "10110111001" => data <= X"001001D4";
         WHEN "10110111010" => data <= X"951DA59C";
         WHEN "10110111011" => data <= X"04D09AE0";
         WHEN "10110111100" => data <= X"2CFCFF07";
         WHEN "10110111101" => data <= X"04C078E0";
         WHEN "10110111110" => data <= X"00F0A018";
         WHEN "10110111111" => data <= X"001001D4";
         WHEN "10111000000" => data <= X"AE1DA59C";
         WHEN "10111000001" => data <= X"04D09AE0";
         WHEN "10111000010" => data <= X"26FCFF07";
         WHEN "10111000011" => data <= X"04C078E0";
         WHEN "10111000100" => data <= X"7CFDFF03";
         WHEN "10111000101" => data <= X"0000001B";
         WHEN "10111000110" => data <= X"01009C9F";
         WHEN "10111000111" => data <= X"00883CE4";
         WHEN "10111001000" => data <= X"B6FFFF13";
         WHEN "10111001001" => data <= X"04D09AE0";
         WHEN "10111001010" => data <= X"F5FFFF03";
         WHEN "10111001011" => data <= X"00F0A018";
         WHEN "10111001100" => data <= X"AFFCFF07";
         WHEN "10111001101" => data <= X"00000015";
         WHEN "10111001110" => data <= X"ADFCFF07";
         WHEN "10111001111" => data <= X"FF004BA7";
         WHEN "10111010000" => data <= X"D0FF5A9F";
         WHEN "10111010001" => data <= X"020020AA";
         WHEN "10111010010" => data <= X"08883AE2";
         WHEN "10111010011" => data <= X"FF004BA6";
         WHEN "10111010100" => data <= X"00D031E2";
         WHEN "10111010101" => data <= X"008831E2";
         WHEN "10111010110" => data <= X"D0FF529E";
         WHEN "10111010111" => data <= X"69FDFF03";
         WHEN "10111011000" => data <= X"008852E2";
         WHEN "10111011001" => data <= X"C91DA59C";
         WHEN "10111011010" => data <= X"0CFEFF03";
         WHEN "10111011011" => data <= X"00008018";
         WHEN "10111011100" => data <= X"1A000010";
         WHEN "10111011101" => data <= X"080020AA";
         WHEN "10111011110" => data <= X"0888D6E2";
         WHEN "10111011111" => data <= X"0100DE9F";
         WHEN "10111100000" => data <= X"040020AA";
         WHEN "10111100001" => data <= X"00883EE4";
         WHEN "10111100010" => data <= X"48000010";
         WHEN "10111100011" => data <= X"00B0DCE2";
         WHEN "10111100100" => data <= X"0C002186";
         WHEN "10111100101" => data <= X"008830E4";
         WHEN "10111100110" => data <= X"17000010";
         WHEN "10111100111" => data <= X"0004201A";
         WHEN "10111101000" => data <= X"FF0720AA";
         WHEN "10111101001" => data <= X"008834E4";
         WHEN "10111101010" => data <= X"0E000010";
         WHEN "10111101011" => data <= X"008854E4";
         WHEN "10111101100" => data <= X"00F0A018";
         WHEN "10111101101" => data <= X"00F08018";
         WHEN "10111101110" => data <= X"00F06018";
         WHEN "10111101111" => data <= X"D71DA59C";
         WHEN "10111110000" => data <= X"B009849C";
         WHEN "10111110001" => data <= X"F7FBFF07";
         WHEN "10111110010" => data <= X"180B639C";
         WHEN "10111110011" => data <= X"010040AA";
         WHEN "10111110100" => data <= X"07000000";
         WHEN "10111110101" => data <= X"000880AA";
         WHEN "10111110110" => data <= X"E9FFFF03";
         WHEN "10111110111" => data <= X"0000C01A";
         WHEN "10111111000" => data <= X"1500000C";
         WHEN "10111111001" => data <= X"020020AA";
         WHEN "10111111010" => data <= X"010040AA";
         WHEN "10111111011" => data <= X"45FDFF03";
         WHEN "10111111100" => data <= X"0000001B";
         WHEN "10111111101" => data <= X"008830E4";
         WHEN "10111111110" => data <= X"0F000010";
         WHEN "10111111111" => data <= X"020020AA";
         WHEN "11000000000" => data <= X"0000201A";
         WHEN "11000000001" => data <= X"008834E4";
         WHEN "11000000010" => data <= X"3EFDFF13";
         WHEN "11000000011" => data <= X"010040AA";
         WHEN "11000000100" => data <= X"00F0A018";
         WHEN "11000000101" => data <= X"00F08018";
         WHEN "11000000110" => data <= X"00F06018";
         WHEN "11000000111" => data <= X"061EA59C";
         WHEN "11000001000" => data <= X"B009849C";
         WHEN "11000001001" => data <= X"DFFBFF07";
         WHEN "11000001010" => data <= X"180B639C";
         WHEN "11000001011" => data <= X"35FDFF03";
         WHEN "11000001100" => data <= X"049092E2";
         WHEN "11000001101" => data <= X"0888D4E3";
         WHEN "11000001110" => data <= X"0000601A";
         WHEN "11000001111" => data <= X"FF3F34A6";
         WHEN "11000010000" => data <= X"009831E4";
         WHEN "11000010001" => data <= X"08000010";
         WHEN "11000010010" => data <= X"00F0A018";
         WHEN "11000010011" => data <= X"00F06018";
         WHEN "11000010100" => data <= X"00F001D4";
         WHEN "11000010101" => data <= X"271EA59C";
         WHEN "11000010110" => data <= X"00008018";
         WHEN "11000010111" => data <= X"D1FBFF07";
         WHEN "11000011000" => data <= X"180B639C";
         WHEN "11000011001" => data <= X"0000201A";
         WHEN "11000011010" => data <= X"00880EE4";
         WHEN "11000011011" => data <= X"11000010";
         WHEN "11000011100" => data <= X"00F030E2";
         WHEN "11000011101" => data <= X"01007672";
         WHEN "11000011110" => data <= X"009811D4";
         WHEN "11000011111" => data <= X"0100949E";
         WHEN "11000100000" => data <= X"00A078E4";
         WHEN "11000100001" => data <= X"09000010";
         WHEN "11000100010" => data <= X"0000C01B";
         WHEN "11000100011" => data <= X"0000201A";
         WHEN "11000100100" => data <= X"00880EE4";
         WHEN "11000100101" => data <= X"03000010";
         WHEN "11000100110" => data <= X"00000015";
         WHEN "11000100111" => data <= X"04A010D4";
         WHEN "11000101000" => data <= X"04A014E3";
         WHEN "11000101001" => data <= X"0000C01B";
         WHEN "11000101010" => data <= X"98FDFF03";
         WHEN "11000101011" => data <= X"FFFF529E";
         WHEN "11000101100" => data <= X"00003186";
         WHEN "11000101101" => data <= X"01003172";
         WHEN "11000101110" => data <= X"008816E4";
         WHEN "11000101111" => data <= X"F0FFFF13";
         WHEN "11000110000" => data <= X"04D0BAE0";
         WHEN "11000110001" => data <= X"00F06018";
         WHEN "11000110010" => data <= X"08B001D4";
         WHEN "11000110011" => data <= X"048801D4";
         WHEN "11000110100" => data <= X"00F001D4";
         WHEN "11000110101" => data <= X"00008018";
         WHEN "11000110110" => data <= X"B2FBFF07";
         WHEN "11000110111" => data <= X"180B639C";
         WHEN "11000111000" => data <= X"E8FFFF03";
         WHEN "11000111001" => data <= X"0100949E";
         WHEN "11000111010" => data <= X"20737562";
         WHEN "11000111011" => data <= X"6F727265";
         WHEN "11000111100" => data <= X"000A2172";
         WHEN "11000111101" => data <= X"61746144";
         WHEN "11000111110" => data <= X"67617020";
         WHEN "11000111111" => data <= X"61662065";
         WHEN "11001000000" => data <= X"0A746C75";
         WHEN "11001000001" => data <= X"70206900";
         WHEN "11001000010" => data <= X"20656761";
         WHEN "11001000011" => data <= X"6C756166";
         WHEN "11001000100" => data <= X"74000A74";
         WHEN "11001000101" => data <= X"0A6B6369";
         WHEN "11001000110" => data <= X"6C6C6100";
         WHEN "11001000111" => data <= X"216E6769";
         WHEN "11001001000" => data <= X"3F3F000A";
         WHEN "11001001001" => data <= X"000A3F3F";
         WHEN "11001001010" => data <= X"676E6970";
         WHEN "11001001011" => data <= X"7464000A";
         WHEN "11001001100" => data <= X"000A626C";
         WHEN "11001001101" => data <= X"626C7469";
         WHEN "11001001110" => data <= X"6152000A";
         WHEN "11001001111" => data <= X"2165676E";
         WHEN "11001010000" => data <= X"7953000A";
         WHEN "11001010001" => data <= X"6C616373";
         WHEN "11001010010" => data <= X"54000A6C";
         WHEN "11001010011" => data <= X"21706172";
         WHEN "11001010100" => data <= X"7242000A";
         WHEN "11001010101" => data <= X"0A6B6165";
         WHEN "11001010110" => data <= X"65684300";
         WHEN "11001010111" => data <= X"6E696B63";
         WHEN "11001011000" => data <= X"616C2067";
         WHEN "11001011001" => data <= X"70207473";
         WHEN "11001011010" => data <= X"20656761";
         WHEN "11001011011" => data <= X"6620666F";
         WHEN "11001011100" => data <= X"6873616C";
         WHEN "11001011101" => data <= X"706D6520";
         WHEN "11001011110" => data <= X"000A7974";
         WHEN "11001011111" => data <= X"73616C46";
         WHEN "11001100000" => data <= X"72652068";
         WHEN "11001100001" => data <= X"21726F72";
         WHEN "11001100010" => data <= X"7245000A";
         WHEN "11001100011" => data <= X"6E697361";
         WHEN "11001100100" => data <= X"616C2067";
         WHEN "11001100101" => data <= X"70207473";
         WHEN "11001100110" => data <= X"20656761";
         WHEN "11001100111" => data <= X"4620666F";
         WHEN "11001101000" => data <= X"6873616C";
         WHEN "11001101001" => data <= X"7257000A";
         WHEN "11001101010" => data <= X"6E697469";
         WHEN "11001101011" => data <= X"65742067";
         WHEN "11001101100" => data <= X"73207473";
         WHEN "11001101101" => data <= X"65757165";
         WHEN "11001101110" => data <= X"2065636E";
         WHEN "11001101111" => data <= X"66206F74";
         WHEN "11001110000" => data <= X"6873616C";
         WHEN "11001110001" => data <= X"56000A2E";
         WHEN "11001110010" => data <= X"66697265";
         WHEN "11001110011" => data <= X"676E6979";
         WHEN "11001110100" => data <= X"73657420";
         WHEN "11001110101" => data <= X"65732074";
         WHEN "11001110110" => data <= X"6E657571";
         WHEN "11001110111" => data <= X"66206563";
         WHEN "11001111000" => data <= X"206D6F72";
         WHEN "11001111001" => data <= X"73616C66";
         WHEN "11001111010" => data <= X"000A2E68";
         WHEN "11001111011" => data <= X"74736554";
         WHEN "11001111100" => data <= X"69616620";
         WHEN "11001111101" => data <= X"3A64656C";
         WHEN "11001111110" => data <= X"20642520";
         WHEN "11001111111" => data <= X"7830203A";
         WHEN "11010000000" => data <= X"2F205825";
         WHEN "11010000001" => data <= X"7830203D";
         WHEN "11010000010" => data <= X"000A5825";
         WHEN "11010000011" => data <= X"73616C46";
         WHEN "11010000100" => data <= X"65742068";
         WHEN "11010000101" => data <= X"6F207473";
         WHEN "11010000110" => data <= X"2E79616B";
         WHEN "11010000111" => data <= X"43000A0A";
         WHEN "11010001000" => data <= X"37342D53";
         WHEN "11010001001" => data <= X"79532033";
         WHEN "11010001010" => data <= X"6D657473";
         WHEN "11010001011" => data <= X"6F727020";
         WHEN "11010001100" => data <= X"6D617267";
         WHEN "11010001101" => data <= X"676E696D";
         WHEN "11010001110" => data <= X"726F6620";
         WHEN "11010001111" => data <= X"73797320";
         WHEN "11010010000" => data <= X"736D6574";
         WHEN "11010010001" => data <= X"206E6F20";
         WHEN "11010010010" => data <= X"70696863";
         WHEN "11010010011" => data <= X"704F000A";
         WHEN "11010010100" => data <= X"69726E65";
         WHEN "11010010101" => data <= X"62206373";
         WHEN "11010010110" => data <= X"64657361";
         WHEN "11010010111" => data <= X"72697620";
         WHEN "11010011000" => data <= X"6C617574";
         WHEN "11010011001" => data <= X"6F725020";
         WHEN "11010011010" => data <= X"79746F74";
         WHEN "11010011011" => data <= X"0A2E6570";
         WHEN "11010011100" => data <= X"69754200";
         WHEN "11010011101" => data <= X"7620646C";
         WHEN "11010011110" => data <= X"69737265";
         WHEN "11010011111" => data <= X"203A6E6F";
         WHEN "11010100000" => data <= X"30206153";
         WHEN "11010100001" => data <= X"65462033";
         WHEN "11010100010" => data <= X"30322062";
         WHEN "11010100011" => data <= X"31203432";
         WHEN "11010100100" => data <= X"39353A31";
         WHEN "11010100101" => data <= X"2036323A";
         WHEN "11010100110" => data <= X"0A544543";
         WHEN "11010100111" => data <= X"2049000A";
         WHEN "11010101000" => data <= X"43206D61";
         WHEN "11010101001" => data <= X"25205550";
         WHEN "11010101010" => data <= X"666F2064";
         WHEN "11010101011" => data <= X"20642520";
         WHEN "11010101100" => data <= X"6E6E7572";
         WHEN "11010101101" => data <= X"20676E69";
         WHEN "11010101110" => data <= X"00207461";
         WHEN "11010101111" => data <= X"64256425";
         WHEN "11010110000" => data <= X"2564252E";
         WHEN "11010110001" => data <= X"484D2064";
         WHEN "11010110010" => data <= X"0A0A2E7A";
         WHEN "11010110011" => data <= X"776F4400";
         WHEN "11010110100" => data <= X"616F6C6E";
         WHEN "11010110101" => data <= X"64203A64";
         WHEN "11010110110" => data <= X"0A656E6F";
         WHEN "11010110111" => data <= X"61655200";
         WHEN "11010111000" => data <= X"676E6964";
         WHEN "11010111001" => data <= X"646F6320";
         WHEN "11010111010" => data <= X"61742065";
         WHEN "11010111011" => data <= X"0A656C62";
         WHEN "11010111100" => data <= X"776F4400";
         WHEN "11010111101" => data <= X"616F6C6E";
         WHEN "11010111110" => data <= X"73203A64";
         WHEN "11010111111" => data <= X"61207465";
         WHEN "11011000000" => data <= X"65726464";
         WHEN "11011000001" => data <= X"3D207373";
         WHEN "11011000010" => data <= X"25783020";
         WHEN "11011000011" => data <= X"45000A58";
         WHEN "11011000100" => data <= X"726F7272";
         WHEN "11011000101" => data <= X"6F6E202C";
         WHEN "11011000110" => data <= X"6F727020";
         WHEN "11011000111" => data <= X"6D617267";
         WHEN "11011001000" => data <= X"616F6C20";
         WHEN "11011001001" => data <= X"21646564";
         WHEN "11011001010" => data <= X"754A000A";
         WHEN "11011001011" => data <= X"6E69706D";
         WHEN "11011001100" => data <= X"6F742067";
         WHEN "11011001101" => data <= X"6F727020";
         WHEN "11011001110" => data <= X"6D617267";
         WHEN "11011001111" => data <= X"45000A6D";
         WHEN "11011010000" => data <= X"726F7272";
         WHEN "11011010001" => data <= X"6F6E202C";
         WHEN "11011010010" => data <= X"6F727020";
         WHEN "11011010011" => data <= X"6D617267";
         WHEN "11011010100" => data <= X"206E6920";
         WHEN "11011010101" => data <= X"73616C46";
         WHEN "11011010110" => data <= X"000A2168";
         WHEN "11011010111" => data <= X"74746553";
         WHEN "11011011000" => data <= X"20676E69";
         WHEN "11011011001" => data <= X"676F7270";
         WHEN "11011011010" => data <= X"6F6D202E";
         WHEN "11011011011" => data <= X"000A6564";
         WHEN "11011011100" => data <= X"74746553";
         WHEN "11011011101" => data <= X"20676E69";
         WHEN "11011011110" => data <= X"69726576";
         WHEN "11011011111" => data <= X"6D202E66";
         WHEN "11011100000" => data <= X"0A65646F";
         WHEN "11011100001" => data <= X"206F4E00";
         WHEN "11011100010" => data <= X"676F7270";
         WHEN "11011100011" => data <= X"206D6172";
         WHEN "11011100100" => data <= X"73657270";
         WHEN "11011100101" => data <= X"0A746E65";
         WHEN "11011100110" => data <= X"6F725000";
         WHEN "11011100111" => data <= X"6D617267";
         WHEN "11011101000" => data <= X"206E6920";
         WHEN "11011101001" => data <= X"206D656D";
         WHEN "11011101010" => data <= X"6D6F7266";
         WHEN "11011101011" => data <= X"25783020";
         WHEN "11011101100" => data <= X"6F742058";
         WHEN "11011101101" => data <= X"25783020";
         WHEN "11011101110" => data <= X"53000A58";
         WHEN "11011101111" => data <= X"63746977";
         WHEN "11011110000" => data <= X"20646568";
         WHEN "11011110001" => data <= X"73206F74";
         WHEN "11011110010" => data <= X"2D74666F";
         WHEN "11011110011" => data <= X"736F6962";
         WHEN "11011110100" => data <= X"7753000A";
         WHEN "11011110101" => data <= X"68637469";
         WHEN "11011110110" => data <= X"74206465";
         WHEN "11011110111" => data <= X"6C46206F";
         WHEN "11011111000" => data <= X"0A687361";
         WHEN "11011111001" => data <= X"69775300";
         WHEN "11011111010" => data <= X"65686374";
         WHEN "11011111011" => data <= X"6F742064";
         WHEN "11011111100" => data <= X"52445320";
         WHEN "11011111101" => data <= X"000A6D61";
         WHEN "11011111110" => data <= X"61656C50";
         WHEN "11011111111" => data <= X"63206573";
         WHEN "11100000000" => data <= X"676E6168";
         WHEN "11100000001" => data <= X"6F742065";
         WHEN "11100000010" => data <= X"65687420";
         WHEN "11100000011" => data <= X"52445320";
         WHEN "11100000100" => data <= X"62204D41";
         WHEN "11100000101" => data <= X"742A2079";
         WHEN "11100000110" => data <= X"6F4E000A";
         WHEN "11100000111" => data <= X"6F727020";
         WHEN "11100001000" => data <= X"6D617267";
         WHEN "11100001001" => data <= X"616F6C20";
         WHEN "11100001010" => data <= X"20646564";
         WHEN "11100001011" => data <= X"53206E69";
         WHEN "11100001100" => data <= X"6D615244";
         WHEN "11100001101" => data <= X"50000A21";
         WHEN "11100001110" => data <= X"72676F72";
         WHEN "11100001111" => data <= X"64206D61";
         WHEN "11100010000" => data <= X"2073656F";
         WHEN "11100010001" => data <= X"20746F6E";
         WHEN "11100010010" => data <= X"20746966";
         WHEN "11100010011" => data <= X"46206E69";
         WHEN "11100010100" => data <= X"6873616C";
         WHEN "11100010101" => data <= X"43000A21";
         WHEN "11100010110" => data <= X"61706D6F";
         WHEN "11100010111" => data <= X"65206572";
         WHEN "11100011000" => data <= X"726F7272";
         WHEN "11100011001" => data <= X"20746120";
         WHEN "11100011010" => data <= X"58257830";
         WHEN "11100011011" => data <= X"30203A20";
         WHEN "11100011100" => data <= X"20582578";
         WHEN "11100011101" => data <= X"30203D21";
         WHEN "11100011110" => data <= X"0A582578";
         WHEN "11100011111" => data <= X"6D6F4300";
         WHEN "11100100000" => data <= X"65726170";
         WHEN "11100100001" => data <= X"6E6F6420";
         WHEN "11100100010" => data <= X"43000A65";
         WHEN "11100100011" => data <= X"6B636568";
         WHEN "11100100100" => data <= X"20676E69";
         WHEN "11100100101" => data <= X"74206669";
         WHEN "11100100110" => data <= X"66206568";
         WHEN "11100100111" => data <= X"6873616C";
         WHEN "11100101000" => data <= X"20736920";
         WHEN "11100101001" => data <= X"74706D65";
         WHEN "11100101010" => data <= X"2E2E2E79";
         WHEN "11100101011" => data <= X"7453000A";
         WHEN "11100101100" => data <= X"20747261";
         WHEN "11100101101" => data <= X"73616C66";
         WHEN "11100101110" => data <= X"72652068";
         WHEN "11100101111" => data <= X"20657361";
         WHEN "11100110000" => data <= X"6C637963";
         WHEN "11100110001" => data <= X"6F662065";
         WHEN "11100110010" => data <= X"61702072";
         WHEN "11100110011" => data <= X"30206567";
         WHEN "11100110100" => data <= X"0A582578";
         WHEN "11100110101" => data <= X"61745300";
         WHEN "11100110110" => data <= X"70207472";
         WHEN "11100110111" => data <= X"72676F72";
         WHEN "11100111000" => data <= X"696D6D61";
         WHEN "11100111001" => data <= X"6620676E";
         WHEN "11100111010" => data <= X"6873616C";
         WHEN "11100111011" => data <= X"7250000A";
         WHEN "11100111100" => data <= X"6172676F";
         WHEN "11100111101" => data <= X"6E696D6D";
         WHEN "11100111110" => data <= X"69662067";
         WHEN "11100111111" => data <= X"6873696E";
         WHEN "11101000000" => data <= X"000A6465";
         WHEN "11101000001" => data <= X"63656843";
         WHEN "11101000010" => data <= X"676E696B";
         WHEN "11101000011" => data <= X"20666920";
         WHEN "11101000100" => data <= X"73616C66";
         WHEN "11101000101" => data <= X"73692068";
         WHEN "11101000110" => data <= X"69642720";
         WHEN "11101000111" => data <= X"27797472";
         WHEN "11101001000" => data <= X"6C46000A";
         WHEN "11101001001" => data <= X"20687361";
         WHEN "11101001010" => data <= X"65207369";
         WHEN "11101001011" => data <= X"7974706D";
         WHEN "11101001100" => data <= X"72652820";
         WHEN "11101001101" => data <= X"64657361";
         WHEN "11101001110" => data <= X"0A0A2E29";
         WHEN "11101001111" => data <= X"61745300";
         WHEN "11101010000" => data <= X"6E697472";
         WHEN "11101010001" => data <= X"69732067";
         WHEN "11101010010" => data <= X"656C706D";
         WHEN "11101010011" => data <= X"52445320";
         WHEN "11101010100" => data <= X"6D206D61";
         WHEN "11101010101" => data <= X"68636D65";
         WHEN "11101010110" => data <= X"2E6B6365";
         WHEN "11101010111" => data <= X"57000A0A";
         WHEN "11101011000" => data <= X"69746972";
         WHEN "11101011001" => data <= X"2E2E676E";
         WHEN "11101011010" => data <= X"56000A2E";
         WHEN "11101011011" => data <= X"66697265";
         WHEN "11101011100" => data <= X"676E6979";
         WHEN "11101011101" => data <= X"0A2E2E2E";
         WHEN "11101011110" => data <= X"72724500";
         WHEN "11101011111" => data <= X"4020726F";
         WHEN "11101100000" => data <= X"58257830";
         WHEN "11101100001" => data <= X"30203A20";
         WHEN "11101100010" => data <= X"20582578";
         WHEN "11101100011" => data <= X"30203D21";
         WHEN "11101100100" => data <= X"0A582578";
         WHEN "11101100101" => data <= X"20724E00";
         WHEN "11101100110" => data <= X"6520666F";
         WHEN "11101100111" => data <= X"726F7272";
         WHEN "11101101000" => data <= X"6F662073";
         WHEN "11101101001" => data <= X"20646E75";
         WHEN "11101101010" => data <= X"6425203A";
         WHEN "11101101011" => data <= X"654D000A";
         WHEN "11101101100" => data <= X"6568636D";
         WHEN "11101101101" => data <= X"64206B63";
         WHEN "11101101110" => data <= X"2C656E6F";
         WHEN "11101101111" => data <= X"20642520";
         WHEN "11101110000" => data <= X"6F727265";
         WHEN "11101110001" => data <= X"0A0A7372";
         WHEN "11101110010" => data <= X"6B6E5500";
         WHEN "11101110011" => data <= X"6E776F6E";
         WHEN "11101110100" => data <= X"646F6320";
         WHEN "11101110101" => data <= X"50002165";
         WHEN "11101110110" => data <= X"72676F72";
         WHEN "11101110111" => data <= X"74206D61";
         WHEN "11101111000" => data <= X"62206F6F";
         WHEN "11101111001" => data <= X"74206769";
         WHEN "11101111010" => data <= X"6966206F";
         WHEN "11101111011" => data <= X"6E692074";
         WHEN "11101111100" => data <= X"666F5320";
         WHEN "11101111101" => data <= X"6F696274";
         WHEN "11101111110" => data <= X"61202C73";
         WHEN "11101111111" => data <= X"74726F62";
         WHEN "11110000000" => data <= X"21676E69";
         WHEN "11110000001" => data <= X"6143000A";
         WHEN "11110000010" => data <= X"746F6E6E";
         WHEN "11110000011" => data <= X"6F727020";
         WHEN "11110000100" => data <= X"6D617267";
         WHEN "11110000101" => data <= X"616C6620";
         WHEN "11110000110" => data <= X"202C6873";
         WHEN "11110000111" => data <= X"726F6261";
         WHEN "11110001000" => data <= X"676E6974";
         WHEN "11110001001" => data <= X"44000A21";
         WHEN "11110001010" => data <= X"6C6E776F";
         WHEN "11110001011" => data <= X"3A64616F";
         WHEN "11110001100" => data <= X"20746120";
         WHEN "11110001101" => data <= X"58257830";
         WHEN "11110001110" => data <= X"6556000A";
         WHEN "11110001111" => data <= X"69666972";
         WHEN "11110010000" => data <= X"69746163";
         WHEN "11110010001" => data <= X"65206E6F";
         WHEN "11110010010" => data <= X"726F7272";
         WHEN "11110010011" => data <= X"20746120";
         WHEN "11110010100" => data <= X"58257830";
         WHEN "11110010101" => data <= X"30203A20";
         WHEN "11110010110" => data <= X"20582578";
         WHEN "11110010111" => data <= X"30203D21";
         WHEN "11110011000" => data <= X"0A582578";
         WHEN "11110011010" => data <= X"EFBEADDE";
         WHEN "11110011011" => data <= X"01000000";
         WHEN "11110011100" => data <= X"02000000";
         WHEN "11110011101" => data <= X"03000000";
         WHEN "11110011110" => data <= X"04000000";
         WHEN "11110011111" => data <= X"05000000";
         WHEN "11110100000" => data <= X"06000000";
         WHEN "11110100001" => data <= X"07000000";
         WHEN OTHERS => data <= X"00000000";
      END CASE;
   END PROCESS TheRom;

END platform_independent;
